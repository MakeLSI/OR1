# dff1_r
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Tue Jun 16 07:57:59 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO dff1_r
    CLASS core ;
    FOREIGN dff1_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 59.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 2.0 14.0 4.0 16.0 ;
        END
    END CK
    PIN Q
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 57.0 4.5 58.0 20.5 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT 18.0 9.0 20.0 11.0 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 59.5 30.0 ;
        RECT 1.0 20.5 3.0 30.0 ;
        RECT 10.5 20.5 12.5 30.0 ;
        RECT 17.0 20.5 19.0 30.0 ;
        RECT 27.0 20.5 29.0 30.0 ;
        RECT 33.5 20.5 35.5 30.0 ;
        RECT 43.5 20.5 45.5 30.0 ;
        RECT 53.0 20.5 55.0 30.0 ;
	END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 59.5 1.0 ;
        RECT 1.0 -1.0 3.0 4.5 ;
        RECT 10.5 -1.0 12.5 4.5 ;
        RECT 17.0 -1.0 19.0 4.5 ;
        RECT 27.0 -1.0 29.0 4.5 ;
        RECT 33.5 -1.0 35.5 4.5 ;
        RECT 43.5 -1.0 45.5 4.5 ;
        RECT 53.5 -1.0 55.5 4.5 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        RECT 23.0 12.5 34.5 13.5 ;
        RECT 39.5 4.5 40.5 6.5 ;
        RECT 28.0 6.0 32.5 7.0 ;
        RECT 25.0 15.5 37.5 16.5 ;
        RECT 14.5 4.5 15.5 10.0 ;
        RECT 14.0 15.5 23.0 16.5 ;
        RECT 9.5 18.5 11.5 19.5 ;
        RECT 23.0 18.5 28.0 19.5 ;        
        RECT 32.0 18.5 32.5 19.5 ;
        RECT 40.5 18.5 44.5 19.5 ;
        RECT 48.5 8.5 51.0 9.5 ;
        RECT 51.0 6.0 54.0 7.0 ;
        RECT 52.0 18.5 54.0 19.5 ;
        RECT 18.0 9.0 20.0 11.0 ;
        RECT 2.0 14.0 4.0 16.0 ;
        RECT 51.0 18.5 52.0 20.5 ;
        RECT 54.5 8.0 55.5 17.5 ;
        RECT 51.0 4.5 52.0 6.0 ;
        RECT 47.5 4.5 48.5 20.5 ;
        RECT 5.0 4.5 6.0 20.5 ;
        RECT 36.5 12.5 39.5 13.5 ;
        RECT 18.0 12.5 21.0 13.5 ;
        RECT 40.5 5.5 44.5 6.5 ;
        RECT 30.5 4.5 31.5 6.0 ;
        RECT 24.0 2.5 25 10.5 ;
        RECT 15.5 6.0 21.0 7.0 ;
        RECT 14.0 9.0 15.0 15.5 ;
        RECT 14.5 16.5 15.5 20.5 ;
        RECT 9.5 12.5 11.0 13.5 ;
        RECT 8.5 4.5 9.5 20.5 ;
        RECT 23.0 19.5 24.0 20.5 ;
        RECT 31.0 18.5 32.0 20.5 ;
        RECT 39.5 18.5 40.5 20.5 ;
        RECT 48.5 16.0 51.0 17.0 ;
        RECT 44.5 13.5 47.5 14.5 ;
        RECT 25.0 9.5 28.5 10.5 ;
        RECT 9.5 6.0 11.5 7.0 ;
        RECT 43.5 20.5 45.5 30.0 ;
        RECT 27.0 20.5 29.0 30.0 ;
        RECT 10.5 20.5 12.5 30.0 ;
        RECT 1.0 20.5 3.0 30.0 ;
        RECT 22.0 2.5 25.0 4.5 ;
        RECT 57.0 4.5 58.0 20.5 ;
        RECT 17.0 20.5 19.0 30.0 ;
        RECT 33.5 20.5 35.5 30.0 ;
        RECT 53.0 20.5 55.0 30.0 ;

        LAYER ML1 ;
      # VIA 5 23.5 dcont
        RECT 4.0 22.5 6 24.5 ;
      # VIA 2 25.5 dcont
        RECT 1.0 24.5 3 26.5 ;
      # VIA 5 25.5 dcont
        RECT 4.0 24.5 6 26.5 ;
      # VIA 2 23.5 dcont
        RECT 1.0 22.5 3 24.5 ;
      # VIA 2 3.5 dcont
        RECT 1.0 2.5 3 4.5 ;
      # VIA 5 3.5 dcont
        RECT 4 2.5 6 4.5 ;
      # VIA 2 21.5 dcont
        RECT 1 20.5 3 22.5 ;
      # VIA 5 21.5 dcont
        RECT 4 20.5 6 22.5 ;
      # VIA 3 15 pcont
        RECT 2 14 4 16 ;
      # VIA 54 3.5 dcont
        RECT 53 2.5 55 4.5 ;
      # VIA 14.5 25.5 dcont
        RECT 13.5 24.5 15.5 26.5 ;
      # VIA 55 7 pcont
        RECT 54 6 56 8 ;
      # VIA 39.5 3.5 dcont
        RECT 38.5 2.5 40.5 4.5 ;
      # VIA 14.5 23.5 dcont
        RECT 13.5 22.5 15.5 24.5 ;
      # VIA 23 25.5 dcont
        RECT 22 24.5 24 26.5 ;
      # VIA 14.5 3.5 dcont
        RECT 13.5 2.5 15.5 4.5 ;
      # VIA 40.5 13.5 pcont
        RECT 39.5 12.5 41.5 14.5 ;
      # VIA 45.5 18.5 pcont
        RECT 44.5 17.5 46.5 19.5 ;
      # VIA 29.5 10 pcont
        RECT 28.5 9 30.5 11 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 12.5 18.5 pcont
        RECT 11.5 17.5 13.5 19.5 ;
      # VIA 34.5 25.5 dcont
        RECT 33.5 24.5 35.5 26.5 ;
      # VIA 22 13 pcont
        RECT 21 12 23 14 ;
      # VIA 18 23.5 dcont
        RECT 17 22.5 19 24.5 ;
      # VIA 45.5 6.5 pcont
        RECT 44.5 5.5 46.5 7.5 ;
      # VIA 23 23.5 dcont
        RECT 22 22.5 24 24.5 ;
      # VIA 54 25.5 dcont
        RECT 53 24.5 55 26.5 ;
      # VIA 27 6.5 pcont
        RECT 26 5.5 28 7.5 ;
      # VIA 39.5 25.5 dcont
        RECT 38.5 24.5 40.5 26.5 ;
      # VIA 34.5 21.5 dcont
        RECT 33.5 20.5 35.5 22.5 ;
      # VIA 44.5 25.5 dcont
        RECT 43.5 24.5 45.5 26.5 ;
      # VIA 28 23.5 dcont
        RECT 27 22.5 29 24.5 ;
      # VIA 11.5 23.5 dcont
        RECT 10.5 22.5 12.5 24.5 ;
      # VIA 8.5 3.5 dcont
        RECT 7.5 2.5 9.5 4.5 ;
      # VIA 28 21.5 dcont
        RECT 27 20.5 29 22.5 ;
      # VIA 23 3.5 dcont
        RECT 22 2.5 24 4.5 ;
      # VIA 28 3.5 dcont
        RECT 27 2.5 29 4.5 ;
      # VIA 44.5 3.5 dcont
        RECT 43.5 2.5 45.5 4.5 ;
      # VIA 11.5 3.5 dcont
        RECT 10.5 2.5 12.5 4.5 ;
      # VIA 22 6.5 pcont
        RECT 21 5.5 23 7.5 ;
      # VIA 43.5 14 pcont
        RECT 42.5 13 44.5 15 ;
      # VIA 14.5 21.5 dcont
        RECT 13.5 20.5 15.5 22.5 ;
      # VIA 34.5 23.5 dcont
        RECT 33.5 22.5 35.5 24.5 ;
      # VIA 33.5 6.5 pcont
        RECT 32.5 5.5 34.5 7.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 34.5 3.5 dcont
        RECT 33.5 2.5 35.5 4.5 ;
      # VIA 47.5 23.5 dcont
        RECT 46.5 22.5 48.5 24.5 ;
      # VIA 31 21.5 dcont
        RECT 30 20.5 32 22.5 ;
      # VIA 39.5 21.5 dcont
        RECT 38.5 20.5 40.5 22.5 ;
      # VIA 24 16 pcont
        RECT 23 15 25 17 ;
      # VIA 44.5 21.5 dcont
        RECT 43.5 20.5 45.5 22.5 ;
      # VIA 18 3.5 dcont
        RECT 17 2.5 19 4.5 ;
      # VIA 18 25.5 dcont
        RECT 17 24.5 19 26.5 ;
      # VIA 57 25.5 dcont
        RECT 56 24.5 58 26.5 ;
      # VIA 29 18.5 pcont
        RECT 28 17.5 30 19.5 ;
      # VIA 57 21.5 dcont
        RECT 56 20.5 58 22.5 ;
      # VIA 28 25.5 dcont
        RECT 27 24.5 29 26.5 ;
      # VIA 23 21.5 dcont
        RECT 22 20.5 24 22.5 ;
      # VIA 38.5 16.5 pcont
        RECT 37.5 15.5 39.5 17.5 ;
      # VIA 52 9 pcont
        RECT 51 8 53 10 ;
      # VIA 17 13 pcont
        RECT 16 12 18 14 ;
      # VIA 31 3.5 dcont
        RECT 30 2.5 32 4.5 ;
      # VIA 18 21.5 dcont
        RECT 17 20.5 19 22.5 ;
      # VIA 31 25.5 dcont
        RECT 30 24.5 32 26.5 ;
      # VIA 52 16.5 pcont
        RECT 51 15.5 53 17.5 ;
      # VIA 19 10 pcont
        RECT 18 9 20 11 ;
      # VIA 8.5 21.5 dcont
        RECT 7.5 20.5 9.5 22.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 11.5 25.5 dcont
        RECT 10.5 24.5 12.5 26.5 ;
      # VIA 57 3.5 dcont
        RECT 56 2.5 58 4.5 ;
      # VIA 54 23.5 dcont
        RECT 53 22.5 55 24.5 ;
      # VIA 35.5 13 pcont
        RECT 34.5 12 36.5 14 ;
      # VIA 47.5 21.5 dcont
        RECT 46.5 20.5 48.5 22.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 39.5 23.5 dcont
        RECT 38.5 22.5 40.5 24.5 ;
      # VIA 54 21.5 dcont
        RECT 53 20.5 55 22.5 ;
      # VIA 44.5 23.5 dcont
        RECT 43.5 22.5 45.5 24.5 ;
      # VIA 31 23.5 dcont
        RECT 30 22.5 32 24.5 ;
      # VIA 8.5 23.5 dcont
        RECT 7.5 22.5 9.5 24.5 ;
      # VIA 57 23.5 dcont
        RECT 56 22.5 58 24.5 ;
      # VIA 12 13 pcont
        RECT 11 12 13 14 ;
      # VIA 11.5 21.5 dcont
        RECT 10.5 20.5 12.5 22.5 ;
      # VIA 55 18.5 pcont
        RECT 54 17.5 56 19.5 ;
      # VIA 47.5 3.5 dcont
        RECT 46.5 2.5 48.5 4.5 ;
      # VIA 33.5 18.5 pcont
        RECT 32.5 17.5 34.5 19.5 ;
      # VIA 8.5 25.5 dcont
        RECT 7.5 24.5 9.5 26.5 ;
      # VIA 12.5 6.5 pcont
        RECT 11.5 5.5 13.5 7.5 ;
      # VIA 47.5 25.5 dcont
        RECT 46.5 24.5 48.5 26.5 ;
      # VIA 6.5 15.5 pcont
        RECT 5.5 14.5 7.5 16.5 ;
	END
END dff1_r

END LIBRARY
