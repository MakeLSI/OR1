# OR1_stdcells.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run & Edited by akita11, 200603

version 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;
MANUFACTURINGGRID 0.1 ;

LAYER ML1
 TYPE		ROUTING ;
 DIRECTION	HORIZONTAL ;
 PITCH		3 ;
 OFFSET	1 ;
 WIDTH		1 ;
 SPACING	1 ;
 RESISTANCE	RPERSQ 0.07 ;
 CAPACITANCE	CPERSQDIST 3e-05 ;
END ML1

LAYER VIA1
 TYPE	CUT ;
 SPACING	1.0 ;
END VIA1

LAYER ML2
 TYPE		ROUTING ;
 DIRECTION	VERTICAL ;
 PITCH		3 ;
 OFFSET	1 ;
 WIDTH		1 ;
 SPACING	1 ;
 RESISTANCE	RPERSQ 0.07 ;
 CAPACITANCE	CPERSQDIST 1.7e-05 ;
END ML2

LAYER VIA2
 TYPE	CUT ;
 SPACING	1.0 ;
END VIA2

LAYER ML3
 TYPE		ROUTING ;
 DIRECTION	HORIZONTAL ;
 PITCH		3 ;
 OFFSET	1 ;
 WIDTH		1 ;
 SPACING	1 ;
 RESISTANCE	RPERSQ 0.07 ;
 CAPACITANCE	CPERSQDIST 7e-06 ;
END ML3

LAYER DM_VIA1
 TYPE	CUT ;
 SPACING	1.0 ;
END DM_VIA1

LAYER DM_VIA2
 TYPE	CUT ;
 SPACING	1.0 ;
END DM_VIA2

VIA M2_M1 DEFAULT
 LAYER ML1 ;
  RECT -1.0 -1.0 1.0 1.0 ;
 LAYER VIA1 ;
  RECT -0.5 -0.5 0.5 0.5 ;
 LAYER ML2 ;
  RECT -1.0 -1.0 1.0 1.0 ;
 LAYER DM_VIA1 ;
  RECT -1.0 -1.0 1.0 1.0 ;
END M2_M1

VIA M3_M2 DEFAULT
 LAYER ML2 ;
  RECT -1.0 -1.0 1.0 1.0 ;
 LAYER VIA2 ;
  RECT -0.5 -0.5 0.5 0.5 ;
 LAYER ML3 ;
  RECT -1.0 -1.0 1.0 1.0 ;
 LAYER DM_VIA2 ;
  RECT -1.0 -1.0 1.0 1.0 ;
END M3_M2

#MACRO dcont
# CLASS CORE ;
# SIZE 2.0 BY 2.0 ;
# ORIGIN 0.0 0.0 ;
# OBS
# END
#END dcont
#MACRO pcont
# CLASS CORE ;
# SIZE 2.0 BY 2.0 ;
# ORIGIN 0.0 0.0 ;
# OBS
# END
#END pcont

MACRO VIA1
 CLASS CORE ;
 SIZE 2.0 BY 2.0 ;
 ORIGIN 0.0 0.0 ;
 OBS
 END
END VIA1

VIARULE viagen21 GENERATE
 LAYER ML1 ;
  DIRECTION HORIZONTAL ;
  WIDTH 1.0 TO 60 ;
  OVERHANG 0.5 ;
  METALOVERHANG 0 ;
 LAYER ML2 ;
  DIRECTION VERTICAL ;
  WIDTH 1.0 TO 60 ;
  OVERHANG 0.5 ;
  METALOVERHANG 0 ;
 LAYER VIA1 ;
  RECT -0.5 -0.5 0.5 0.5 ;
  SPACING 1 BY 1 ;
END viagen21

VIARULE viagen32 GENERATE
 LAYER ML3 ;
  DIRECTION HORIZONTAL ;
  WIDTH 1.0 TO 60 ;
  OVERHANG 0.5 ;
  METALOVERHANG 0 ;
 LAYER ML2 ;
  DIRECTION VERTICAL ;
  WIDTH 1.0 TO 60 ;
  OVERHANG 0.5 ;
  METALOVERHANG 0 ;
 LAYER VIA2 ;
  RECT -0.5 -0.5 0.5 0.5 ;
  SPACING 1 BY 1 ;
END viagen32

VIARULE TURN1 GENERATE
 LAYER ML1 ;
  DIRECTION HORIZONTAL ;
 LAYER ML1 ;
  DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
 LAYER ML2 ;
  DIRECTION HORIZONTAL ;
 LAYER ML2 ;
  DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
 LAYER ML3 ;
  DIRECTION HORIZONTAL ;
 LAYER ML3 ;
  DIRECTION VERTICAL ;
END TURN3

MACRO FILL
 CLASS CORE ;
 FOREIGN FILL 0.0 0.0 ;
 ORIGIN 0.0 0.0 ;
 SIZE 3.0 BY 29.0 ;
 SYMMETRY X ;
 SITE core ;
 PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
  PORT
   LAYER ML1 ;
    RECT -0.5 -1.0 3.5 1.0 ;
  END
 END VSS
 PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
  PORT
   LAYER ML1 ;
    RECT -0.5 28.0 3.5 30.0 ;
  END
 END VDD
END FILL

MACRO an21
    CLASS core ;
    FOREIGN an21 0.0 0.0;
    ORIGIN 0.0 0.0 ;
    SYMMETRY X Y ;
    SIZE 12.5 BY 29.0 ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 12.5 12.0 14.5 ;
        LAYER ML1 ;
        RECT 10.0 12.5 12.0 14.5 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 12.5 6.0 14.5 ;
        LAYER ML1 ;
        RECT 4.0 12.5 6.0 14.5 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 10.0 3.0 12.0 ;
        LAYER ML1 ;
        RECT 1.0 10.0 3.0 12.0 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 6.5 9.5 6.5 9.5 3.5 ;
        WIDTH 2 ;
        PATH 6.5 0.0 6.5 3.5 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 18.0 7.5 18.0 7.5 8.5 1.5 8.5 1.5 3.5 ;
        WIDTH 2 ;
        PATH 7.5 21.5 7.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        LAYER ML1 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 8 10.5 pcont
        RECT 7 9.5 9 11.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 6.5 3.5 dcont
        RECT 5.5 2.5 7.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 9.5 3.5 dcont
        RECT 8.5 2.5 10.5 4.5 ;
    END
END an21
MACRO an31
    CLASS core ;
    FOREIGN an31 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    SYMMETRY X Y ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.0 12.5 15.0 14.5 ;
        LAYER ML1 ;
        RECT 13.0 12.5 15.0 14.5 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 12.5 6.0 14.5 ;
        LAYER ML1 ;
        RECT 4.0 12.5 6.0 14.5 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 9.5 3.0 11.5 ;
        LAYER ML1 ;
        RECT 1.0 9.5 3.0 11.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 9.5 9.0 11.5 ;
        LAYER ML1 ;
        RECT 7.0 9.5 9.0 11.5 ;
        END
    END C
    OBS
        LAYER ML1 ;
        WIDTH 1 ;
        PATH 13.5 25.5 13.5 4.0 11.5 4.0 11.5 3.8 ;
        WIDTH 1.4 ;
        PATH 13.5 22.3 13.5 25.5 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 10.5 21.5 10.5 28.5 ;
        WIDTH 2 ;
        PATH 8.5 0.0 8.5 3.5 ;
        WIDTH 1.4 ;
        PATH 7.5 22.3 7.5 25.5 ;
        WIDTH 1 ;
        PATH 7.5 21.5 7.5 18.0 ;
        
        WIDTH 1 ;
        PATH 1.5 21.5 1.5 18.0 10.5 18.0 10.5 8.0 2.0 8.0 2.0 3.8 ;
        WIDTH 2 ;
        PATH 4.5 21.5 4.5 28.5 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        LAYER ML1 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 11.5 3.5 dcont
        RECT 10.5 2.5 12.5 4.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 8.5 3.5 dcont
        RECT 7.5 2.5 9.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 11 10.5 pcont
        RECT 10 9.5 12 11.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
    END
END an31
MACRO an41
    CLASS core ;
    FOREIGN an41 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 18.5 BY 29.0 ;
    SYMMETRY X Y ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 16.0 12.5 18.0 14.5 ;
        LAYER ML1 ;
        RECT 16.0 12.5 18.0 14.5 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 19.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 12.5 6.0 14.5 ;
        LAYER ML1 ;
        RECT 4.0 12.5 6.0 14.5 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 10.0 12.5 12.0 14.5 ;
        LAYER ML1 ;
        RECT 10.0 12.5 12.0 14.5 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 7.0 10.0 9.0 12.0 ;
        LAYER ML2 ;
        RECT 7.0 10.0 9.0 12.0 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 15.5 3.0 17.5 ;
        LAYER ML1 ;
        RECT 1.0 15.5 3.0 17.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 19.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 2 ;
        PATH 10.5 0.0 10.5 3.5 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 2 ;
        PATH 7.5 21.5 7.5 29.0 ;
        WIDTH 1 ;
        PATH 4.5 21.5 4.5 18.0 13.5 18.0 13.5 8.0 1.5 8.0 1.5 3.8 ;
        WIDTH 1 ;
        PATH 10.5 21.5 10.5 18.0 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 13.5 21.5 13.5 28.5 ;
        WIDTH 1.4 ;
        PATH 13.5 22.3 13.5 25.5 ;
        WIDTH 1 ;
        PATH 16.5 21.5 16.5 5.0 14.0 5.0 14.0 3.8 ;
        WIDTH 1.4 ;
        PATH 16.5 22.3 16.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 16.5 21.5 dcont
        RECT 15.5 20.5 17.5 22.5 ;
      # VIA 14 10.5 pcont
        RECT 13 9.5 15 11.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 16.5 25.5 dcont
        RECT 15.5 24.5 17.5 26.5 ;
      # VIA 16.5 23.5 dcont
        RECT 15.5 22.5 17.5 24.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
    END
END an41
MACRO buf1
    CLASS core ;
    FOREIGN buf1 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 9.5 BY 29.0 ;
#    SYMMETRY X ;
    PIN Y
        DIRECTION OUTPUT ;
#        USE SIGNAL ;
        PORT
#        LAYER ML2 ;
#	      RECT 7.0 14.0 9.0 16.0 ;
        LAYER ML1 ;
#              RECT 7.0 14.0 9.0 16.0 ;
              RECT 7.0 3.5 8.0 22.0 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
       	      RECT -0.5 28.0 10.0 30.0 ;
              RECT 3.5 20.5 5.5 29.5 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
              RECT -0.5 -1.0 10.0 1.0 ;
	      RECT 3.5 0.0 5.5 4.5 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
#        USE SIGNAL ;
        PORT
#        LAYER ML2 ;
#              RECT 1.0 14.0 3.0 16.0 ;
        LAYER ML1 ;
              RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
	WIDTH 1.0 ;
	PATH 1.5 21.5 1.5 18.0 4.5 18.0 4.5 7.5 2.0 7.5 2.0 3.8 ;
        RECT 6.5 2.5 8.5 4.5 ;
        RECT 6.5 20.5 8.5 26.5 ;
#	RECT 1.5 3.0 2.5 8.0 ;
#	RECT 1.5 7.0 5.0 8.0 ;
#	RECT 4.0 7.0 5.0 18.5 ;
#	RECT 1.0 17.5 5.0 18.5 ;
#	RECT 1.0 17.5 2.0 22.0 ;
#       RECT 4 10.5 6 12.5 ;
       RECT 0.5 2.5 2.5 4.5 ;
       RECT 0.5 20.5 2.5 26.5 ;
    END
END buf1
MACRO buf2
    CLASS core ;
    FOREIGN buf2 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 14.0 9.0 16.0 ;
        LAYER ML1 ;
        RECT 7.0 14.0 9.0 16.0 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 10.5 21.0 10.5 28.5 ;
        WIDTH 2 ;
        PATH 10.5 1.0 10.5 3.5 ;
        WIDTH 1 ;
        PATH 7.5 3.9 7.5 20.5 ;
        WIDTH 1.4 ;
        PATH 7.5 22.3 7.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.5 ;
        WIDTH 2 ;
        PATH 4.5 21.0 4.5 28.5 ;
        WIDTH 1 ;
        PATH 2.0 20.5 2.0 18.0 4.5 18.0 4.5 7.5 2.0 7.5 2.0 3.8 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 5 11.5 pcont
        RECT 4 10.5 6 12.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
    END
END buf2
MACRO buf4
    CLASS core ;
    FOREIGN buf4 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 18.5 BY 29.0 ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.0 15.0 15.0 17.0 ;
        LAYER ML1 ;
        RECT 13.0 15.0 15.0 17.0 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 19.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 19.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 16.5 1.0 16.5 3.5 ;
        WIDTH 2 ;
        PATH 16.5 21.5 16.5 28.5 ;
        WIDTH 1 ;
        PATH 13.5 3.5 13.5 20.5 ;
        WIDTH 1 ;
        PATH 7.5 8.5 13.5 8.5 ;
        WIDTH 1 ;
        PATH 7.5 7.5 13.5 7.5 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 10.5 21.5 10.5 28.5 ;
        WIDTH 2 ;
        PATH 10.5 1.0 10.5 3.5 ;
        
        
        WIDTH 1 ;
        PATH 7.5 3.5 7.5 20.5 ;
        WIDTH 1.4 ;
        PATH 7.5 21.5 7.5 25.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.5 ;
        WIDTH 2 ;
        PATH 4.5 21.2 4.5 28.5 ;
        WIDTH 1 ;
        PATH 1.5 20.5 1.5 18.0 4.5 18.0 4.5 7.5 2.0 7.5 2.0 3.5 ;
        WIDTH 1.4 ;
        PATH 1.5 21.5 1.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
      # VIA 16.5 23.5 dcont
        RECT 15.5 22.5 17.5 24.5 ;
      # VIA 16.5 25.5 dcont
        RECT 15.5 24.5 17.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 16.5 21.5 dcont
        RECT 15.5 20.5 17.5 22.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
      # VIA 5 11.5 pcont
        RECT 4 10.5 6 12.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 16.5 3.5 dcont
        RECT 15.5 2.5 17.5 4.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
    END
END buf4
MACRO buf8
    CLASS core ;
    FOREIGN buf8 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SYMMETRY X Y  ;
    SIZE 30.5 BY 29.0 ;
        PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 24.0 14.0 26.0 16.0 ;
        LAYER ML1 ;
        RECT 24.0 14.0 26.0 16.0 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 31.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 31.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 2.0 14.0 4.0 16.0 ;
        LAYER ML1 ;
        RECT 2.0 14.0 4.0 16.0 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 28.5 0.5 28.5 3.5 ;
        WIDTH 2 ;
        PATH 28.5 21.3 28.5 28.5 ;
        WIDTH 1 ;
        PATH 25.5 3.9 25.5 20.5 ;
        WIDTH 1.4 ;
        PATH 25.5 22.3 25.5 25.5 ;
        WIDTH 2 ;
        PATH 22.5 0.5 22.5 3.5 ;
        WIDTH 2 ;
        PATH 22.5 21.5 22.5 28.5 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 19.5 3.9 19.5 20.5 ;
        WIDTH 1.4 ;
        PATH 19.5 21.5 19.5 25.5 ;
        WIDTH 1 ;
        PATH 7.5 8.5 25.5 8.5 ;
        WIDTH 1 ;
        PATH 7.5 7.5 25.5 7.5 ;
        WIDTH 2 ;
        PATH 16.5 0.5 16.5 3.5 ;
        WIDTH 2 ;
        PATH 16.5 21.6 16.5 28.5 ;
        
        
        WIDTH 1 ;
        PATH 13.5 3.9 13.5 20.5 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 10.5 21.5 10.5 28.5 ;
        WIDTH 2 ;
        PATH 10.5 0.5 10.5 3.5 ;
        WIDTH 1 ;
        PATH 7.5 4.0 7.5 20.5 ;
        WIDTH 1.4 ;
        PATH 7.5 21.5 7.5 25.5 ;
        WIDTH 2 ;
        PATH 4.5 0.5 4.5 3.5 ;
        WIDTH 2 ;
        PATH 4.5 21.5 4.5 28.5 ;
        WIDTH 1 ;
        PATH 2.0 20.5 2.0 18.0 4.5 18.0 4.5 7.5 2.0 7.5 2.0 3.5 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1.4 ;
        PATH 13.5 21.5 13.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
      # VIA 25.5 25.5 dcont
        RECT 24.5 24.5 26.5 26.5 ;
      # VIA 28.5 25.5 dcont
        RECT 27.5 24.5 29.5 26.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 16.5 23.5 dcont
        RECT 15.5 22.5 17.5 24.5 ;
      # VIA 16.5 25.5 dcont
        RECT 15.5 24.5 17.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 28.5 3.5 dcont
        RECT 27.5 2.5 29.5 4.5 ;
      # VIA 5 11.5 pcont
        RECT 4 10.5 6 12.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 19.5 25.5 dcont
        RECT 18.5 24.5 20.5 26.5 ;
      # VIA 16.5 21.5 dcont
        RECT 15.5 20.5 17.5 22.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
      # VIA 25.5 23.5 dcont
        RECT 24.5 22.5 26.5 24.5 ;
      # VIA 19.5 23.5 dcont
        RECT 18.5 22.5 20.5 24.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 28.5 21.5 dcont
        RECT 27.5 20.5 29.5 22.5 ;
      # VIA 16.5 3.5 dcont
        RECT 15.5 2.5 17.5 4.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 25.5 3.5 dcont
        RECT 24.5 2.5 26.5 4.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 19.5 3.5 dcont
        RECT 18.5 2.5 20.5 4.5 ;
      # VIA 28.5 23.5 dcont
        RECT 27.5 22.5 29.5 24.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 25.5 21.5 dcont
        RECT 24.5 20.5 26.5 22.5 ;
      # VIA 19.5 21.5 dcont
        RECT 18.5 20.5 20.5 22.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
    END
END buf8
MACRO cinv
    CLASS core ;
    FOREIGN cinv 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 11.5 BY 29.0 ;
    PIN OE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END OE
    PIN YB
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 9.0 7.5 11.0 9.5 ;
        LAYER ML1 ;
        RECT 9.0 7.5 11.0 9.5 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 12.0 30.0 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 6.5 11.5 8.5 13.5 ;
        LAYER ML1 ;
        RECT 6.5 11.5 8.5 13.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 12.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1.4 ;
        PATH 1.5 22.1 1.5 25.5 ;
        WIDTH 1 ;
        PATH 2.0 24.5 2.0 18.0 5.0 18.0 5.0 8.0 2.0 8.0 2.0 3.5 ;
        WIDTH 2 ;
        PATH 4.5 21.5 4.5 28.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.5 ;
        
        
        WIDTH 1.4 ;
        PATH 9.5 22.3 9.5 25.5 ;
        WIDTH 1 ;
        PATH 9.5 20.5 9.5 18.0 10.0 18.0 10.0 8.5 9.5 8.5 9.5 3.5 ;
        
        LAYER ML1 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 9.5 25.5 dcont
        RECT 8.5 24.5 10.5 26.5 ;
      # VIA 5.5 15.5 pcont
        RECT 4.5 14.5 6.5 16.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 9.5 23.5 dcont
        RECT 8.5 22.5 10.5 24.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 9.5 21.5 dcont
        RECT 8.5 20.5 10.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 9.5 3.5 dcont
        RECT 8.5 2.5 10.5 4.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
    END
END cinv
MACRO dff1
    CLASS core ;
    FOREIGN dff1 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 52.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN Q
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.5 51.5 12.5 ;
        LAYER ML1 ;
        RECT 49.5 10.5 51.5 12.5 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 52.5 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 52.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        RECT 15 2.5 18 4.5 ;
        WIDTH 1 ;
        PATH 16.0 3.5 16.0 4.0 17.5 4.0 17.5 9.5 22.0 9.5 ;
        WIDTH 1 ;
        PATH 50.5 3.0 50.5 25.7 ;
        WIDTH 1.4 ;
        PATH 50.0 22.3 50.0 25.5 ;
        WIDTH 1.4 ;
        PATH 50.0 22.3 50.0 25.5 ;
        WIDTH 2 ;
        PATH 47.0 21.5 47.0 28.2 ;
        WIDTH 2 ;
        PATH 47.0 3.5 47.0 1.0 ;
        WIDTH 1 ;
        PATH 44.0 3.5 44.0 6.0 47.5 6.0 47.5 19.0 44.0 19.0 44.0 21.5 ;
        WIDTH 1.4 ;
        PATH 44.0 22.3 44.0 25.5 ;
        WIDTH 1 ;
        PATH 45.0 16.5 41.0 16.5 ;
        WIDTH 1 ;
        PATH 45.0 8.5 41.0 8.5 ;
        WIDTH 1 ;
        PATH 41.0 25.5 41.0 3.4 ;
        WIDTH 1.4 ;
        PATH 40.5 22.3 40.5 25.5 ;
        WIDTH 1 ;
        PATH 36.5 13.5 41.0 13.5 ;
        WIDTH 2 ;
        PATH 37.5 21.5 37.5 28.2 ;
        WIDTH 2 ;
        PATH 37.5 3.5 37.5 1.0 ;
        WIDTH 1 ;
        PATH 32.5 3.5 32.5 6.5 38.5 6.5 ;
        WIDTH 1 ;
        PATH 38.5 19.0 32.5 19.0 32.5 21.5 ;
        WIDTH 1.4 ;
        PATH 32.5 22.3 32.5 25.5 ;
        WIDTH 2 ;
        PATH 27.5 21.5 27.5 28.2 ;
        WIDTH 2 ;
        PATH 27.5 3.5 27.5 1.0 ;
        
        
        WIDTH 1 ;
        PATH 26.5 19.0 24.5 19.0 24.5 21.5 24.0 21.5 ;
        WIDTH 1.4 ;
        PATH 24.0 22.3 24.0 25.5 ;
        WIDTH 1 ;
        PATH 24.0 6.5 24.0 3.4 ;
        WIDTH 1 ;
        PATH 20.0 6.5 26.5 6.5 ;
        WIDTH 1 ;
        PATH 10.0 13.0 33.5 13.0 ;
        WIDTH 2 ;
        PATH 21.0 21.5 21.0 28.2 ;
        WIDTH 2 ;
        PATH 21.0 3.5 21.0 1.0 ;
        WIDTH 1 ;
        PATH 8.0 3.3 8.0 9.0 7.5 9.0 7.5 16.0 31.0 16.0 ;
        WIDTH 1 ;
        PATH 16.0 21.5 16.0 18.5 22.0 18.5 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 14.5 6.5 8.0 6.5 ;
        WIDTH 2 ;
        PATH 11.0 21.5 11.0 28.2 ;
        WIDTH 2 ;
        PATH 11.0 3.5 11.0 1.0 ;
        WIDTH 1 ;
        PATH 8.0 25.5 8.0 16.0 ;
        WIDTH 1.4 ;
        PATH 7.5 22.3 7.5 25.5 ;
        WIDTH 2 ;
        PATH 4.5 21.5 4.5 28.2 ;
        WIDTH 2 ;
        PATH 4.5 3.5 4.5 1.2 ;
        WIDTH 1 ;
        PATH 5.5 6.5 1.5 6.5 ;
        WIDTH 1 ;
        PATH 5.5 18.5 1.5 18.5 ;
        WIDTH 1 ;
        PATH 5.0 13.0 1.5 13.0 ;
        WIDTH 1 ;
        PATH 1.5 3.5 1.5 21.5 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 40.5 25.5 dcont
        RECT 39.5 24.5 41.5 26.5 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 26.5 18.5 pcont
        RECT 25.5 17.5 27.5 19.5 ;
      # VIA 40.5 3.5 dcont
        RECT 39.5 2.5 41.5 4.5 ;
      # VIA 48 18.5 pcont
        RECT 47 17.5 49 19.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 50 23.5 dcont
        RECT 49 22.5 51 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 24 23.5 dcont
        RECT 23 22.5 25 24.5 ;
      # VIA 37.5 23.5 dcont
        RECT 36.5 22.5 38.5 24.5 ;
      # VIA 47 21.5 dcont
        RECT 46 20.5 48 22.5 ;
      # VIA 32.5 23.5 dcont
        RECT 31.5 22.5 33.5 24.5 ;
      # VIA 44 25.5 dcont
        RECT 43 24.5 45 26.5 ;
      # VIA 40.5 21.5 dcont
        RECT 39.5 20.5 41.5 22.5 ;
      # VIA 28.5 13 pcont
        RECT 27.5 12 29.5 14 ;
      # VIA 50 3.5 dcont
        RECT 49 2.5 51 4.5 ;
      # VIA 47 23.5 dcont
        RECT 46 22.5 48 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 44 3.5 dcont
        RECT 43 2.5 45 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 45 16.5 pcont
        RECT 44 15.5 46 17.5 ;
      # VIA 24 25.5 dcont
        RECT 23 24.5 25 26.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 24 3.5 dcont
        RECT 23 2.5 25 4.5 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 45 8.5 pcont
        RECT 44 7.5 46 9.5 ;
      # VIA 31.5 16.5 pcont
        RECT 30.5 15.5 32.5 17.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 50 21.5 dcont
        RECT 49 20.5 51 22.5 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 50 25.5 dcont
        RECT 49 24.5 51 26.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 37.5 21.5 dcont
        RECT 36.5 20.5 38.5 22.5 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 32.5 21.5 dcont
        RECT 31.5 20.5 33.5 22.5 ;
      # VIA 24 21.5 dcont
        RECT 23 20.5 25 22.5 ;
      # VIA 40.5 23.5 dcont
        RECT 39.5 22.5 41.5 24.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 44 23.5 dcont
        RECT 43 22.5 45 24.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 36.5 13.5 pcont
        RECT 35.5 12.5 37.5 14.5 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 37.5 3.5 dcont
        RECT 36.5 2.5 38.5 4.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 37.5 25.5 dcont
        RECT 36.5 24.5 38.5 26.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 32.5 25.5 dcont
        RECT 31.5 24.5 33.5 26.5 ;
      # VIA 20 6.5 pcont
        RECT 19 5.5 21 7.5 ;
      # VIA 47 25.5 dcont
        RECT 46 24.5 48 26.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 38.5 6.5 pcont
        RECT 37.5 5.5 39.5 7.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 15 13 pcont
        RECT 14 12 16 14 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
      # VIA 44 21.5 dcont
        RECT 43 20.5 45 22.5 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 38.5 18.5 pcont
        RECT 37.5 17.5 39.5 19.5 ;
      # VIA 33.5 13.5 pcont
        RECT 32.5 12.5 34.5 14.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 32.5 3.5 dcont
        RECT 31.5 2.5 33.5 4.5 ;
      # VIA 48 6.5 pcont
        RECT 47 5.5 49 7.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 47 3.5 dcont
        RECT 46 2.5 48 4.5 ;
    END
END dff1
MACRO dff1_r
    CLASS core ;
    FOREIGN dff1_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 58.5 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 59.0 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN Q
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 56.0 10.5 58.0 12.5 ;
        LAYER ML1 ;
        RECT 56.0 10.5 58.0 12.5 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 59.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 1.5 21.3 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 5.0 20.5 5.0 3.8 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 8.5 3.5 8.5 21.4 ;
        WIDTH 1 ;
        PATH 11.5 13.0 8.5 13.0 ;
        WIDTH 1 ;
        PATH 12.0 19.0 8.5 19.0 ;
        WIDTH 1 ;
        PATH 12.3 6.5 8.5 6.5 ;
        WIDTH 2 ;
        PATH 11.0 3.6 11.0 1.5 ;
        WIDTH 2 ;
        PATH 11.0 21.8 11.0 28.5 ;
        WIDTH 1.4 ;
        PATH 14.0 22.3 14.0 25.5 ;
        WIDTH 1 ;
        PATH 14.5 25.8 14.5 16.0 ;
        WIDTH 2 ;
        PATH 17.5 3.5 17.5 1.5 ;
        WIDTH 2 ;
        PATH 17.5 21.8 17.5 28.5 ;
        WIDTH 1 ;
        PATH 21.5 6.5 14.5 6.5 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 23.0 21.5 23.0 19.0 28.5 19.0 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 16.0 37.5 16.0 ;
        WIDTH 2 ;
        PATH 27.5 3.5 27.5 1.5 ;
        WIDTH 2 ;
        PATH 27.5 21.8 27.5 28.5 ;
        WIDTH 1 ;
        PATH 16.5 13.0 40.4 13.0 ;
        WIDTH 1 ;
        PATH 26.5 6.5 33.0 6.5 ;
        WIDTH 1 ;
        PATH 30.5 6.5 30.5 3.5 ;
        WIDTH 1.4 ;
        PATH 30.5 22.3 30.5 25.5 ;
        WIDTH 1 ;
        PATH 33.3 19.0 31.0 19.0 31.0 21.8 30.8 21.8 ;
        
        
        WIDTH 2 ;
        PATH 34.0 3.8 34.0 1.5 ;
        WIDTH 2 ;
        PATH 34.0 21.8 34.0 28.5 ;
        WIDTH 1.4 ;
        PATH 39.0 22.3 39.0 25.5 ;
        WIDTH 1 ;
        PATH 45.3 19.0 39.5 19.0 39.5 21.8 ;
        WIDTH 1 ;
        PATH 39.5 3.8 39.5 6.0 44.9 6.0 ;
        WIDTH 2 ;
        PATH 44.0 3.5 44.0 1.2 ;
        WIDTH 2 ;
        PATH 44.0 21.8 44.0 28.5 ;
        WIDTH 1 ;
        PATH 43.0 14.0 47.5 14.0 ;
        WIDTH 1.4 ;
        PATH 47.0 22.3 47.0 25.5 ;
        WIDTH 1 ;
        PATH 47.5 25.8 47.5 3.5 ;
        WIDTH 1 ;
        PATH 51.5 9.0 47.5 9.0 ;
        WIDTH 1 ;
        PATH 51.5 16.5 47.5 16.5 ;
        WIDTH 1.4 ;
        PATH 50.5 22.3 50.5 25.5 ;
        WIDTH 1 ;
        PATH 51.0 3.8 51.0 6.0 54.5 6.0 54.5 19.0 51.0 19.0 51.0 21.8 ;
        WIDTH 2 ;
        PATH 53.5 3.5 53.5 1.5 ;
        WIDTH 2 ;
        PATH 53.5 21.8 53.5 28.5 ;
        WIDTH 1.4 ;
        PATH 56.5 22.3 56.5 25.5 ;
        WIDTH 1.4 ;
        PATH 56.5 22.3 56.5 25.5 ;
        WIDTH 1 ;
        PATH 57.0 3.5 57.0 26.0 ;
        WIDTH 1 ;
        PATH 24.0 4.0 24.0 10.0 29.0 10.0 ;
        RECT 21.5 2.5 24.5 4.5 ;
        
        LAYER ML1 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 53.5 3.5 dcont
        RECT 52.5 2.5 54.5 4.5 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 54.5 7 pcont
        RECT 53.5 6 55.5 8 ;
      # VIA 39 3.5 dcont
        RECT 38 2.5 40 4.5 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 40 13.5 pcont
        RECT 39 12.5 41 14.5 ;
      # VIA 45 18.5 pcont
        RECT 44 17.5 46 19.5 ;
      # VIA 29 10 pcont
        RECT 28 9 30 11 ;
      # VIA 50.5 21.5 dcont
        RECT 49.5 20.5 51.5 22.5 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 34 25.5 dcont
        RECT 33 24.5 35 26.5 ;
      # VIA 21.5 13 pcont
        RECT 20.5 12 22.5 14 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 45 6.5 pcont
        RECT 44 5.5 46 7.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 53.5 25.5 dcont
        RECT 52.5 24.5 54.5 26.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 39 25.5 dcont
        RECT 38 24.5 40 26.5 ;
      # VIA 34 21.5 dcont
        RECT 33 20.5 35 22.5 ;
      # VIA 44 25.5 dcont
        RECT 43 24.5 45 26.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 44 3.5 dcont
        RECT 43 2.5 45 4.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 43 14 pcont
        RECT 42 13 44 15 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 34 23.5 dcont
        RECT 33 22.5 35 24.5 ;
      # VIA 33 6.5 pcont
        RECT 32 5.5 34 7.5 ;
      # VIA 50.5 23.5 dcont
        RECT 49.5 22.5 51.5 24.5 ;
      # VIA 34 3.5 dcont
        RECT 33 2.5 35 4.5 ;
      # VIA 47 23.5 dcont
        RECT 46 22.5 48 24.5 ;
      # VIA 30.5 21.5 dcont
        RECT 29.5 20.5 31.5 22.5 ;
      # VIA 39 21.5 dcont
        RECT 38 20.5 40 22.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 44 21.5 dcont
        RECT 43 20.5 45 22.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 56.5 25.5 dcont
        RECT 55.5 24.5 57.5 26.5 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 56.5 21.5 dcont
        RECT 55.5 20.5 57.5 22.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 38 16.5 pcont
        RECT 37 15.5 39 17.5 ;
      # VIA 51.5 9 pcont
        RECT 50.5 8 52.5 10 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 30.5 3.5 dcont
        RECT 29.5 2.5 31.5 4.5 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 30.5 25.5 dcont
        RECT 29.5 24.5 31.5 26.5 ;
      # VIA 51.5 16.5 pcont
        RECT 50.5 15.5 52.5 17.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 50.5 3.5 dcont
        RECT 49.5 2.5 51.5 4.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 56.5 3.5 dcont
        RECT 55.5 2.5 57.5 4.5 ;
      # VIA 53.5 23.5 dcont
        RECT 52.5 22.5 54.5 24.5 ;
      # VIA 35 13 pcont
        RECT 34 12 36 14 ;
      # VIA 47 21.5 dcont
        RECT 46 20.5 48 22.5 ;
      # VIA 50.5 25.5 dcont
        RECT 49.5 24.5 51.5 26.5 ;
      # VIA 39 23.5 dcont
        RECT 38 22.5 40 24.5 ;
      # VIA 53.5 21.5 dcont
        RECT 52.5 20.5 54.5 22.5 ;
      # VIA 44 23.5 dcont
        RECT 43 22.5 45 24.5 ;
      # VIA 30.5 23.5 dcont
        RECT 29.5 22.5 31.5 24.5 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 56.5 23.5 dcont
        RECT 55.5 22.5 57.5 24.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 54.5 18.5 pcont
        RECT 53.5 17.5 55.5 19.5 ;
      # VIA 47 3.5 dcont
        RECT 46 2.5 48 4.5 ;
      # VIA 33 18.5 pcont
        RECT 32 17.5 34 19.5 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 47 25.5 dcont
        RECT 46 24.5 48 26.5 ;
      # VIA 6 15.5 pcont
        RECT 5 14.5 7 16.5 ;
    END
END dff1_r
MACRO dff1m2
    CLASS core ;
    FOREIGN dff1m2 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 52.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.5 51.5 12.5 ;
        LAYER ML1 ;
        RECT 49.5 10.5 51.5 12.5 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 52.5 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 52.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 50.5 3.3 50.5 26.0 ;
        WIDTH 1.4 ;
        PATH 50.0 22.3 50.0 25.5 ;
        WIDTH 2 ;
        PATH 47.0 22.6 47.0 28.5 ;
        WIDTH 2 ;
        PATH 47.0 1.0 47.0 3.4 ;
        WIDTH 1 ;
        PATH 44.5 26.0 44.5 19.0 48.0 19.0 48.0 6.0 44.5 6.0 44.5 3.6 ;
        WIDTH 1.4 ;
        PATH 44.0 22.3 44.0 25.5 ;
        WIDTH 1 ;
        PATH 45.3 8.5 41.0 8.5 ;
        WIDTH 1 ;
        PATH 45.3 16.5 41.0 16.5 ;
        WIDTH 1 ;
        PATH 41.0 21.5 41.0 3.8 ;
        WIDTH 1 ;
        PATH 36.8 14.0 41.0 14.0 ;
        WIDTH 2 ;
        PATH 37.5 1.0 37.5 3.5 ;
        WIDTH 2 ;
        PATH 37.5 22.6 37.5 28.5 ;
        WIDTH 1 ;
        PATH 33.0 3.8 33.0 6.0 38.5 6.0 ;
        WIDTH 1 ;
        PATH 32.5 22.3 32.5 19.0 38.7 19.0 ;
        WIDTH 1.4 ;
        PATH 32.5 22.3 32.5 25.5 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.5 ;
        WIDTH 2 ;
        PATH 27.5 22.0 27.5 28.5 ;
        
        
        WIDTH 1 ;
        PATH 24.0 21.5 24.5 21.5 24.5 18.4 ;
        WIDTH 1.4 ;
        PATH 24.0 22.3 24.0 25.5 ;
        WIDTH 1 ;
        PATH 34.0 13.0 10.3 13.0 ;
        WIDTH 1 ;
        PATH 19.9 6.5 24.0 6.5 24.0 3.5 ;
        WIDTH 2 ;
        PATH 21.0 1.0 21.0 3.5 ;
        WIDTH 2 ;
        PATH 21.0 22.6 21.0 28.5 ;
        WIDTH 1 ;
        PATH 8.1 16.0 31.8 16.0 ;
        WIDTH 1 ;
        PATH 16.0 3.5 16.0 4.0 17.5 4.0 17.5 10.0 22.4 10.0 ;
        WIDTH 1 ;
        PATH 16.0 22.3 16.0 19.0 22.0 19.0 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 14.8 6.5 8.0 6.5 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.5 ;
        WIDTH 1 ;
        PATH 8.0 3.6 8.0 9.5 7.5 9.5 7.5 16.0 8.0 16.0 8.0 26.0 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.5 ;
        WIDTH 2 ;
        PATH 4.5 22.6 4.5 28.5 ;
        WIDTH 1 ;
        PATH 5.9 6.5 1.8 6.5 ;
        WIDTH 1 ;
        PATH 5.6 18.5 1.5 18.5 ;
        WIDTH 1 ;
        PATH 5.0 13.0 1.8 13.0 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 1.5 26.0 1.5 3.6 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 22.5 18.7 22.5 10.0 ;
        WIDTH 1 ;
        PATH 25.0 18.7 25.0 6.8 ;
        WIDTH 1 ;
        PATH 39.0 18.7 39.0 6.5 ;
        LAYER ML1 ;
      # VIA 28.5 13 pcont
        RECT 27.5 12 29.5 14 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 44 25.5 dcont
        RECT 43 24.5 45 26.5 ;
      # VIA 25 18.5 pcont
        RECT 24 17.5 26 19.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 37.5 21.5 dcont
        RECT 36.5 20.5 38.5 22.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 38.5 18.5 dcont
        RECT 37.5 17.5 39.5 19.5 ;
        LAYER ML2 ;
      # VIA 38.5 18.5 dcont
        RECT 37.5 17.5 39.5 19.5 ;
        LAYER ML1 ;
      # VIA 32.5 21.5 dcont
        RECT 31.5 20.5 33.5 22.5 ;
      # VIA 24 21.5 dcont
        RECT 23 20.5 25 22.5 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 25.5 7 dcont
        RECT 24.5 6 26.5 8 ;
        LAYER ML2 ;
      # VIA 25.5 7 dcont
        RECT 24.5 6 26.5 8 ;
        LAYER ML1 ;
      # VIA 48 6.5 pcont
        RECT 47 5.5 49 7.5 ;
      # VIA 15 13 pcont
        RECT 14 12 16 14 ;
      # VIA 25 18.5 dcont
        RECT 24 17.5 26 19.5 ;
        LAYER ML2 ;
      # VIA 25 18.5 dcont
        RECT 24 17.5 26 19.5 ;
        LAYER ML1 ;
      # VIA 38.5 18.5 pcont
        RECT 37.5 17.5 39.5 19.5 ;
      # VIA 33.5 13.5 pcont
        RECT 32.5 12.5 34.5 14.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 48 18.5 pcont
        RECT 47 17.5 49 19.5 ;
      # VIA 37.5 25.5 dcont
        RECT 36.5 24.5 38.5 26.5 ;
      # VIA 36.5 14 pcont
        RECT 35.5 13 37.5 15 ;
      # VIA 32.5 23.5 dcont
        RECT 31.5 22.5 33.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 24 23.5 dcont
        RECT 23 22.5 25 24.5 ;
      # VIA 44 3.5 dcont
        RECT 43 2.5 45 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 47 25.5 dcont
        RECT 46 24.5 48 26.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 50 25.5 dcont
        RECT 49 24.5 51 26.5 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML2 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML1 ;
      # VIA 38.5 6.5 dcont
        RECT 37.5 5.5 39.5 7.5 ;
        LAYER ML2 ;
      # VIA 38.5 6.5 dcont
        RECT 37.5 5.5 39.5 7.5 ;
        LAYER ML1 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 44 23.5 dcont
        RECT 43 22.5 45 24.5 ;
      # VIA 40.5 3.5 dcont
        RECT 39.5 2.5 41.5 4.5 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 31.5 16.5 pcont
        RECT 30.5 15.5 32.5 17.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 38.5 6.5 pcont
        RECT 37.5 5.5 39.5 7.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 40.5 25.5 dcont
        RECT 39.5 24.5 41.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 32.5 3.5 dcont
        RECT 31.5 2.5 33.5 4.5 ;
      # VIA 20 6.5 pcont
        RECT 19 5.5 21 7.5 ;
      # VIA 50 3.5 dcont
        RECT 49 2.5 51 4.5 ;
      # VIA 32.5 25.5 dcont
        RECT 31.5 24.5 33.5 26.5 ;
      # VIA 47 3.5 dcont
        RECT 46 2.5 48 4.5 ;
      # VIA 50 21.5 dcont
        RECT 49 20.5 51 22.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 37.5 23.5 dcont
        RECT 36.5 22.5 38.5 24.5 ;
      # VIA 50 23.5 dcont
        RECT 49 22.5 51 24.5 ;
      # VIA 25.5 7 pcont
        RECT 24.5 6 26.5 8 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 47 23.5 dcont
        RECT 46 22.5 48 24.5 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML2 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML1 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 44 21.5 dcont
        RECT 43 20.5 45 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 24 25.5 dcont
        RECT 23 24.5 25 26.5 ;
      # VIA 45 8.5 pcont
        RECT 44 7.5 46 9.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 37.5 3.5 dcont
        RECT 36.5 2.5 38.5 4.5 ;
      # VIA 47 21.5 dcont
        RECT 46 20.5 48 22.5 ;
      # VIA 40.5 23.5 dcont
        RECT 39.5 22.5 41.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 24 3.5 dcont
        RECT 23 2.5 25 4.5 ;
      # VIA 40.5 21.5 dcont
        RECT 39.5 20.5 41.5 22.5 ;
      # VIA 45 16.5 pcont
        RECT 44 15.5 46 17.5 ;
    END
END dff1m2
MACRO dff1m2_r
    CLASS core ;
    FOREIGN dff1m2_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 58.5 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 59.0 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 56.0 10.5 58.0 12.5 ;
        LAYER ML1 ;
        RECT 56.0 10.5 58.0 12.5 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 59.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 1 ;
        PATH 8.0 26.0 8.0 3.6 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 11.5 13.0 8.3 13.0 ;
        WIDTH 1 ;
        PATH 12.1 18.5 8.0 18.5 ;
        WIDTH 1 ;
        PATH 12.4 6.5 8.3 6.5 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.5 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 16.0 14.5 16.0 14.5 26.0 ;
        WIDTH 2 ;
        PATH 17.5 1.0 17.5 3.5 ;
        WIDTH 2 ;
        PATH 17.5 22.6 17.5 28.5 ;
        WIDTH 1 ;
        PATH 21.3 6.5 14.5 6.5 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 22.5 22.3 22.5 19.0 28.5 19.0 ;
        WIDTH 1 ;
        PATH 22.5 3.5 22.5 4.0 24.0 4.0 24.0 10.0 28.9 10.0 ;
        WIDTH 1 ;
        PATH 14.6 16.0 38.3 16.0 ;
        WIDTH 2 ;
        PATH 27.5 22.6 27.5 28.5 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.5 ;
        WIDTH 1 ;
        PATH 26.4 6.5 30.5 6.5 30.5 3.5 ;
        WIDTH 1 ;
        PATH 40.5 13.0 16.8 13.0 ;
        WIDTH 1.4 ;
        PATH 30.5 22.3 30.5 25.5 ;
        WIDTH 1 ;
        PATH 30.5 21.5 31.0 21.5 31.0 18.4 ;
        
        
        WIDTH 2 ;
        PATH 34.0 22.0 34.0 28.5 ;
        WIDTH 2 ;
        PATH 34.0 1.0 34.0 3.5 ;
        WIDTH 1.4 ;
        PATH 39.0 22.3 39.0 25.5 ;
        WIDTH 1 ;
        PATH 39.0 22.3 39.0 19.0 45.2 19.0 ;
        WIDTH 1 ;
        PATH 39.5 3.8 39.5 6.0 45.0 6.0 ;
        WIDTH 2 ;
        PATH 44.0 22.6 44.0 28.5 ;
        WIDTH 2 ;
        PATH 44.0 1.0 44.0 3.5 ;
        WIDTH 1 ;
        PATH 43.3 14.0 47.5 14.0 ;
        WIDTH 1 ;
        PATH 47.5 21.5 47.5 3.8 ;
        WIDTH 1 ;
        PATH 51.8 16.5 47.5 16.5 ;
        WIDTH 1 ;
        PATH 51.8 8.5 47.5 8.5 ;
        WIDTH 1.4 ;
        PATH 50.5 22.3 50.5 25.5 ;
        WIDTH 1 ;
        PATH 51.0 26.0 51.0 19.0 54.5 19.0 54.5 6.0 51.0 6.0 51.0 3.6 ;
        WIDTH 2 ;
        PATH 53.5 1.0 53.5 3.4 ;
        WIDTH 2 ;
        PATH 53.5 22.6 53.5 28.5 ;
        WIDTH 1.4 ;
        PATH 56.5 22.3 56.5 25.5 ;
        WIDTH 1 ;
        PATH 57.0 3.3 57.0 26.0 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 45.5 18.7 45.5 6.5 ;
        WIDTH 1 ;
        PATH 31.5 18.7 31.5 6.8 ;
        WIDTH 1 ;
        PATH 29.0 18.7 29.0 10.0 ;
        LAYER ML1 ;
      # VIA 5.5 13 pcont
        RECT 4.5 12 6.5 14 ;
      # VIA 35 13 pcont
        RECT 34 12 36 14 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 34 21.5 dcont
        RECT 33 20.5 35 22.5 ;
      # VIA 34 23.5 dcont
        RECT 33 22.5 35 24.5 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 50.5 25.5 dcont
        RECT 49.5 24.5 51.5 26.5 ;
      # VIA 31.5 18.5 pcont
        RECT 30.5 17.5 32.5 19.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 44 21.5 dcont
        RECT 43 20.5 45 22.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 45 18.5 dcont
        RECT 44 17.5 46 19.5 ;
        LAYER ML2 ;
      # VIA 45 18.5 dcont
        RECT 44 17.5 46 19.5 ;
        LAYER ML1 ;
      # VIA 39 21.5 dcont
        RECT 38 20.5 40 22.5 ;
      # VIA 30.5 21.5 dcont
        RECT 29.5 20.5 31.5 22.5 ;
      # VIA 28.5 10 pcont
        RECT 27.5 9 29.5 11 ;
      # VIA 32 7 dcont
        RECT 31 6 33 8 ;
        LAYER ML2 ;
      # VIA 32 7 dcont
        RECT 31 6 33 8 ;
        LAYER ML1 ;
      # VIA 54.5 6.5 pcont
        RECT 53.5 5.5 55.5 7.5 ;
      # VIA 21.5 13 pcont
        RECT 20.5 12 22.5 14 ;
      # VIA 31.5 18.5 dcont
        RECT 30.5 17.5 32.5 19.5 ;
        LAYER ML2 ;
      # VIA 31.5 18.5 dcont
        RECT 30.5 17.5 32.5 19.5 ;
        LAYER ML1 ;
      # VIA 45 18.5 pcont
        RECT 44 17.5 46 19.5 ;
      # VIA 40 13.5 pcont
        RECT 39 12.5 41 14.5 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 54.5 18.5 pcont
        RECT 53.5 17.5 55.5 19.5 ;
      # VIA 44 25.5 dcont
        RECT 43 24.5 45 26.5 ;
      # VIA 43 14 pcont
        RECT 42 13 44 15 ;
      # VIA 39 23.5 dcont
        RECT 38 22.5 40 24.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 30.5 23.5 dcont
        RECT 29.5 22.5 31.5 24.5 ;
      # VIA 50.5 3.5 dcont
        RECT 49.5 2.5 51.5 4.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 53.5 25.5 dcont
        RECT 52.5 24.5 54.5 26.5 ;
      # VIA 34 25.5 dcont
        RECT 33 24.5 35 26.5 ;
      # VIA 56.5 25.5 dcont
        RECT 55.5 24.5 57.5 26.5 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML2 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML1 ;
      # VIA 45 6.5 dcont
        RECT 44 5.5 46 7.5 ;
        LAYER ML2 ;
      # VIA 45 6.5 dcont
        RECT 44 5.5 46 7.5 ;
        LAYER ML1 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 50.5 23.5 dcont
        RECT 49.5 22.5 51.5 24.5 ;
      # VIA 47 3.5 dcont
        RECT 46 2.5 48 4.5 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 38 16.5 pcont
        RECT 37 15.5 39 17.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 45 6.5 pcont
        RECT 44 5.5 46 7.5 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 47 25.5 dcont
        RECT 46 24.5 48 26.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 39 3.5 dcont
        RECT 38 2.5 40 4.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 56.5 3.5 dcont
        RECT 55.5 2.5 57.5 4.5 ;
      # VIA 39 25.5 dcont
        RECT 38 24.5 40 26.5 ;
      # VIA 53.5 3.5 dcont
        RECT 52.5 2.5 54.5 4.5 ;
      # VIA 56.5 21.5 dcont
        RECT 55.5 20.5 57.5 22.5 ;
      # VIA 34 3.5 dcont
        RECT 33 2.5 35 4.5 ;
      # VIA 44 23.5 dcont
        RECT 43 22.5 45 24.5 ;
      # VIA 56.5 23.5 dcont
        RECT 55.5 22.5 57.5 24.5 ;
      # VIA 32 7 pcont
        RECT 31 6 33 8 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 53.5 23.5 dcont
        RECT 52.5 22.5 54.5 24.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 50.5 21.5 dcont
        RECT 49.5 20.5 51.5 22.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML2 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML1 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 30.5 25.5 dcont
        RECT 29.5 24.5 31.5 26.5 ;
      # VIA 51.5 8.5 pcont
        RECT 50.5 7.5 52.5 9.5 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 44 3.5 dcont
        RECT 43 2.5 45 4.5 ;
      # VIA 53.5 21.5 dcont
        RECT 52.5 20.5 54.5 22.5 ;
      # VIA 47 23.5 dcont
        RECT 46 22.5 48 24.5 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 30.5 3.5 dcont
        RECT 29.5 2.5 31.5 4.5 ;
      # VIA 47 21.5 dcont
        RECT 46 20.5 48 22.5 ;
      # VIA 51.5 16.5 pcont
        RECT 50.5 15.5 52.5 17.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
    END
END dff1m2_r
MACRO exnr
    CLASS core ;
    FOREIGN exnr 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 21.0 BY 29.0 ;
        PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 2.0 12.0 5.0 14.0 ;
        LAYER ML1 ;
        RECT 3.0 12.0 5.0 14.0 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 21.5 30.0 ;
        END
    END VDD
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 18.0 12.0 20.0 14.0 ;
        LAYER ML1 ;
        RECT 18.0 12.0 20.0 14.0 ;
        END
    END YB
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 21.5 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 6.0 14.0 8.0 16.0 ;
        LAYER ML1 ;
        RECT 6.0 14.0 8.0 16.0 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 19.0 21.6 19.0 28.5 ;
        WIDTH 1 ;
        PATH 16.5 21.4 16.5 17.5 19.5 17.5 19.5 3.5 ;
        WIDTH 1.4 ;
        PATH 16.0 25.5 16.0 21.5 ;
        WIDTH 1 ;
        PATH 15.5 3.5 15.5 6.0 10.5 6.0 10.5 3.5 ;
        WIDTH 2 ;
        PATH 13.0 1.0 13.0 3.5 ;
        WIDTH 2 ;
        PATH 11.0 21.5 11.0 28.5 ;
        WIDTH 1 ;
        PATH 7.1 14.5 14.5 14.5 ;
        
        
        WIDTH 1 ;
        PATH 1.5 9.0 16.8 9.0 ;
        WIDTH 2 ;
        PATH 7.5 21.8 7.5 28.5 ;
        WIDTH 1 ;
        PATH 4.0 11.5 11.4 11.5 ;
        WIDTH 2 ;
        PATH 6.5 1.0 6.5 3.5 ;
        WIDTH 1 ;
        PATH 4.0 25.5 4.0 19.0 1.5 19.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 11.5 11.5 pcont
        RECT 10.5 10.5 12.5 12.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 19 21.5 dcont
        RECT 18 20.5 20 22.5 ;
      # VIA 19 25.5 dcont
        RECT 18 24.5 20 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 17 9 pcont
        RECT 16 8 18 10 ;
      # VIA 19 23.5 dcont
        RECT 18 22.5 20 24.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 10 3.5 dcont
        RECT 9 2.5 11 4.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 6.5 3.5 dcont
        RECT 5.5 2.5 7.5 4.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 19 3.5 dcont
        RECT 18 2.5 20 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 14.5 14.5 pcont
        RECT 13.5 13.5 15.5 15.5 ;
      # VIA 13 3.5 dcont
        RECT 12 2.5 14 4.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
    END
END exnr
MACRO exor
    CLASS core ;
    FOREIGN exor 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SYMMETRY X Y  ;
    SIZE 21.0 BY 29.0 ;
        PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 18.0 12.0 20.0 14.0 ;
        LAYER ML1 ;
        RECT 18.0 12.0 20.0 14.0 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 3.0 10.0 5.0 12.0 ;
        LAYER ML1 ;
        RECT 3.0 10.0 5.0 12.0 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 21.5 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 21.5 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 6.0 14.0 8.0 16.0 ;
        LAYER ML1 ;
        RECT 6.0 14.0 8.0 16.0 ;
        END
    END A
    OBS
        LAYER ML1 ;
        WIDTH 1.4 ;
        PATH 19.0 21.5 19.0 25.5 ;
        WIDTH 2 ;
        PATH 18.0 1.0 18.0 3.5 ;
        WIDTH 1 ;
        PATH 19.0 21.8 19.0 6.0 15.5 6.0 15.5 3.5 ;
        WIDTH 1 ;
        PATH 16.0 25.5 16.0 18.5 10.0 18.5 10.0 24.8 ;
        WIDTH 2 ;
        PATH 13.0 21.5 13.0 28.5 ;
        WIDTH 1 ;
        PATH 7.0 14.5 14.2 14.5 ;
        WIDTH 2 ;
        PATH 10.0 1.0 10.0 3.5 ;
        WIDTH 1 ;
        PATH 4.0 11.0 11.0 11.0 ;
        WIDTH 2 ;
        PATH 6.5 21.5 6.5 28.5 ;
        WIDTH 1 ;
        PATH 4.5 8.5 4.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 16.7 8.5 1.5 8.5 1.5 25.5 ;
        LAYER ML1 ;
      # VIA 11 11 pcont
        RECT 10 10 12 12 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 19 23.5 dcont
        RECT 18 22.5 20 24.5 ;
      # VIA 19 21.5 dcont
        RECT 18 20.5 20 22.5 ;
      # VIA 6.5 21.5 dcont
        RECT 5.5 20.5 7.5 22.5 ;
      # VIA 13 21.5 dcont
        RECT 12 20.5 14 22.5 ;
      # VIA 10 23.5 dcont
        RECT 9 22.5 11 24.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 10 21.5 dcont
        RECT 9 20.5 11 22.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 16.5 8.5 pcont
        RECT 15.5 7.5 17.5 9.5 ;
      # VIA 18 3.5 dcont
        RECT 17 2.5 19 4.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 10 25.5 dcont
        RECT 9 24.5 11 26.5 ;
      # VIA 15 3.5 dcont
        RECT 14 2.5 16 4.5 ;
      # VIA 6.5 25.5 dcont
        RECT 5.5 24.5 7.5 26.5 ;
      # VIA 10 3.5 dcont
        RECT 9 2.5 11 4.5 ;
      # VIA 6.5 23.5 dcont
        RECT 5.5 22.5 7.5 24.5 ;
      # VIA 19 25.5 dcont
        RECT 18 24.5 20 26.5 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 13 23.5 dcont
        RECT 12 22.5 14 24.5 ;
      # VIA 14 14.5 pcont
        RECT 13 13.5 15 15.5 ;
      # VIA 13 25.5 dcont
        RECT 12 24.5 14 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
    END
END exor
MACRO inv1
    CLASS core ;
    FOREIGN inv1 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
#    SYMMETRY XY ;
    SIZE 6.5 BY 29.0 ;
    SITE core ;
    PIN YB
        DIRECTION OUTPUT ;
        PORT
        LAYER ML1 ;
	      RECT 4.0 3.0 5.0 21.0 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
              RECT -0.5 28.0 7.0 30.0 ;
              RECT 0.5 20.5 2.5 29.5 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
              RECT -0.5 -1.0 7.0 1.0 ;
              RECT 0.5 0.0 2.5 4.5 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
#        LAYER ML2 ;
#	      RECT 1.0 14.0 3.0 16.0 ;
        LAYER ML1 ;
              RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
	LAYER ML1 ;
              RECT 3.5 2.5 5.5 4.5 ;
              RECT 3.5 20.5 5.5 26.5 ;
    END
END inv1
MACRO inv2
    CLASS core ;
    FOREIGN inv2 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 9.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.0 6.0 13.0 ;
        LAYER ML1 ;
        RECT 4.0 11.0 6.0 13.0 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 10.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 10.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
        WIDTH 2 ;
        PATH 7.5 1.0 7.5 3.5 ;
        WIDTH 2 ;
        PATH 7.5 21.5 7.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        LAYER ML1 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
    END
END inv2
MACRO inv4
    CLASS core ;
    FOREIGN inv4 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 10.0 12.0 12.0 ;
        LAYER ML1 ;
        RECT 10.0 10.0 12.0 12.0 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 13.5 0.5 13.5 3.5 ;
        WIDTH 2 ;
        PATH 13.5 21.6 13.5 28.5 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 3.8 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 7.5 0.5 7.5 3.5 ;
        WIDTH 2 ;
        PATH 7.5 21.3 7.5 28.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.3 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 0.5 1.5 3.5 ;
        
        LAYER ML1 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
    END
END inv4
MACRO inv8
    CLASS core ;
    FOREIGN inv8 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 27.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 22.0 10.5 24.0 12.5 ;
        LAYER ML1 ;
        RECT 22.0 10.5 24.0 12.5 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 28.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 28.0 1.0 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.8 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.5 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 2 ;
        PATH 7.5 1.0 7.5 3.8 ;
        WIDTH 2 ;
        PATH 7.5 21.3 7.5 28.5 ;
        WIDTH 1 ;
        PATH 10.5 21.5 10.5 3.5 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 13.5 21.3 13.5 28.5 ;
        WIDTH 1 ;
        PATH 4.8 11.0 22.8 11.0 ;
        WIDTH 2 ;
        PATH 13.5 1.0 13.5 3.8 ;
        WIDTH 1 ;
        PATH 16.5 21.5 16.5 3.5 ;
        WIDTH 1.4 ;
        PATH 19.5 22.3 19.5 25.5 ;
        WIDTH 2 ;
        PATH 19.5 21.3 19.5 28.5 ;
        WIDTH 2 ;
        PATH 19.5 1.0 19.5 3.8 ;
        WIDTH 1 ;
        PATH 22.5 21.5 22.5 3.5 ;
        WIDTH 1.4 ;
        PATH 25.5 22.3 25.5 25.5 ;
        WIDTH 2 ;
        PATH 25.5 21.5 25.5 28.5 ;
        WIDTH 2 ;
        PATH 25.5 1.0 25.5 3.8 ;
        
        LAYER ML1 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 25.5 25.5 dcont
        RECT 24.5 24.5 26.5 26.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 19.5 25.5 dcont
        RECT 18.5 24.5 20.5 26.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 19.5 3.5 dcont
        RECT 18.5 2.5 20.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 25.5 3.5 dcont
        RECT 24.5 2.5 26.5 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 16.5 3.5 dcont
        RECT 15.5 2.5 17.5 4.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 25.5 21.5 dcont
        RECT 24.5 20.5 26.5 22.5 ;
      # VIA 19.5 21.5 dcont
        RECT 18.5 20.5 20.5 22.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
      # VIA 16.5 25.5 dcont
        RECT 15.5 24.5 17.5 26.5 ;
      # VIA 19.5 23.5 dcont
        RECT 18.5 22.5 20.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 16.5 23.5 dcont
        RECT 15.5 22.5 17.5 24.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 16.5 21.5 dcont
        RECT 15.5 20.5 17.5 22.5 ;
      # VIA 25.5 23.5 dcont
        RECT 24.5 22.5 26.5 24.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
    END
END inv8
MACRO na21
    CLASS core ;
    FOREIGN na21 0.0 0.0 ;
#    SYMMETRY X ;
    ORIGIN 0.0 0.0 ;
    SIZE 9.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
#              RECT 6.0 12.0 8.0 14.0 ;
#	       WIDTH 1.0 ;
#	       PATH 5.0 20.5 5.0 18.0 7.5 18.0 7.5 6.5 6.5 6.5 6.5 3.5 ;
	      RECT 6.0 3.0 7.0 7.0 ;
	      RECT 7.0 6.0 8.0 18.5 ;
	      RECT 4.5 17.5 8.0 18.5 ;
	      RECT 4.5 17.5 5.5 21.0 ;
        END
    END YB
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
              RECT 4.0 8.5 6.0 10.5 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
              RECT -0.5 28.0 10.0 30.0 ;
              RECT 0.5 20.5 2.5 29.5 ;
              RECT 6.5 20.5 8.5 29.5 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
              RECT 2.0 14.5 4.0 16.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
              RECT -0.5 -1.0 10.0 1.0 ;
	      RECT 0.5 0.0 2.5 4.5 ;
        END
    END VSS
    OBS
	LAYER ML1 ;
             RECT 3.5 20.5 5.5 26.5 ;
             RECT 5.5 2.5 7.5 4.5 ;
    END
END na21
MACRO na212
    CLASS core ;
    FOREIGN na212 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 8.5 12.0 10.5 ;
        LAYER ML1 ;
        RECT 10.0 8.5 12.0 10.5 ;
        END
    END YB
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 7.0 12.0 9.0 14.0 ;
        LAYER ML2 ;
        RECT 7.0 12.0 9.0 14.0 ;
        END
    END B0
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 10.5 21.5 10.5 28.5 ;
        WIDTH 1 ;
        PATH 7.5 20.5 7.5 18.0 10.5 18.0 10.5 3.5 ;
        WIDTH 1.4 ;
        PATH 7.5 22.3 7.5 25.5 ;
        
        
        WIDTH 1 ;
        PATH 7.5 3.5 7.5 8.0 1.5 8.0 1.5 3.5 ;
        WIDTH 1 ;
        PATH 4.5 1.0 4.5 3.5 ;
        WIDTH 2 ;
        PATH 2.5 21.5 2.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 2.5 25.5 dcont
        RECT 1.5 24.5 3.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 2.5 23.5 dcont
        RECT 1.5 22.5 3.5 24.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 2.5 21.5 dcont
        RECT 1.5 20.5 3.5 22.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
    END
END na212
MACRO na222
    CLASS core ;
    FOREIGN na222 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.0 10.5 15.0 12.5 ;
        LAYER ML1 ;
        RECT 13.0 10.5 15.0 12.5 ;
        END
    END YB
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 10.0 6.0 12.0 ;
        LAYER ML1 ;
        RECT 4.0 10.0 6.0 12.0 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 14.5 12.0 16.5 ;
        LAYER ML1 ;
        RECT 10.0 14.5 12.0 16.5 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 11.5 9.0 13.5 ;
        LAYER ML1 ;
        RECT 7.0 11.5 9.0 13.5 ;
        END
    END B1
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 12.5 21.5 12.5 28.5 ;
        WIDTH 1 ;
        PATH 7.5 20.5 7.5 18.0 13.5 18.0 13.5 8.0 10.5 8.0 10.5 5.5 ;
        WIDTH 1.4 ;
        PATH 7.5 21.5 7.5 25.5 ;
        WIDTH 1 ;
        PATH 13.5 5.5 13.5 2.5 7.5 2.5 7.5 8.0 1.5 8.0 1.5 5.0 ;
        
        
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 5.0 ;
        WIDTH 2 ;
        PATH 2.5 21.5 2.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 13.5 5 dcont
        RECT 12.5 4 14.5 6 ;
      # VIA 12.5 23.5 dcont
        RECT 11.5 22.5 13.5 24.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 2.5 25.5 dcont
        RECT 1.5 24.5 3.5 26.5 ;
      # VIA 12.5 21.5 dcont
        RECT 11.5 20.5 13.5 22.5 ;
      # VIA 2.5 23.5 dcont
        RECT 1.5 22.5 3.5 24.5 ;
      # VIA 10.5 5 dcont
        RECT 9.5 4 11.5 6 ;
      # VIA 4.5 5 dcont
        RECT 3.5 4 5.5 6 ;
      # VIA 2.5 21.5 dcont
        RECT 1.5 20.5 3.5 22.5 ;
      # VIA 12.5 25.5 dcont
        RECT 11.5 24.5 13.5 26.5 ;
      # VIA 7.5 5 dcont
        RECT 6.5 4 8.5 6 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 1.5 5 dcont
        RECT 0.5 4 2.5 6 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
    END
END na222
MACRO na31
    CLASS core ;
    FOREIGN na31 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 12.0 12.0 14.0 ;
        LAYER ML1 ;
        RECT 10.0 12.0 12.0 14.0 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 8.0 9.0 10.0 ;
        LAYER ML1 ;
        RECT 7.0 8.0 9.0 10.0 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 18.0 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 18.0 10.5 18.0 10.5 6.5 9.0 6.5 9.0 3.8 ;
        WIDTH 2 ;
        PATH 7.5 21.6 7.5 28.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 8.5 3.5 dcont
        RECT 7.5 2.5 9.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
        LAYER ML1 ;
        
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 18.0 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 18.0 10.5 18.0 10.5 6.5 9.0 6.5 9.0 3.8 ;
        WIDTH 2 ;
        PATH 7.5 21.6 7.5 28.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 8.5 3.5 dcont
        RECT 7.5 2.5 9.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
    END
END na31
MACRO na41
    CLASS core ;
    FOREIGN na41 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.0 9.5 15.0 11.5 ;
        LAYER ML1 ;
        RECT 13.0 9.5 15.0 11.5 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 12.5 6.0 14.5 ;
        LAYER ML1 ;
        RECT 4.0 12.5 6.0 14.5 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 10.0 6.5 12.0 8.5 ;
        LAYER ML1 ;
        RECT 10.0 6.5 12.0 8.5 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 9.5 9.0 11.5 ;
        LAYER ML1 ;
        RECT 7.0 9.5 9.0 11.5 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 15.5 3.0 17.5 ;
        LAYER ML1 ;
        RECT 1.0 15.5 3.0 17.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 7.5 21.5 7.5 28.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 18.0 13.5 18.0 13.5 4.0 10.6 4.0 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 18.0 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        WIDTH 2 ;
        PATH 13.5 21.5 13.5 28.5 ;
        WIDTH 1.4 ;
        PATH 13.5 22.3 13.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 13.5 25.5 dcont
        RECT 12.5 24.5 14.5 26.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 13.5 21.5 dcont
        RECT 12.5 20.5 14.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
      # VIA 13.5 23.5 dcont
        RECT 12.5 22.5 14.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
    END
END na41
MACRO nr21
    CLASS core ;
    FOREIGN nr21 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 9.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 8.5 9.0 10.5 ;
        LAYER ML1 ;
        RECT 7.0 8.5 9.0 10.5 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 10.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 10.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 4.5 3.5 4.5 6.5 7.5 6.5 7.5 15.5 7.0 15.5 7.0 20.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 7.0 21.5 7.0 25.5 ;
        
        
        WIDTH 2 ;
        PATH 2.0 22.0 2.0 28.5 ;
        WIDTH 2 ;
        PATH 7.5 1.0 7.5 3.5 ;
        
        LAYER ML1 ;
      # VIA 7 21.5 dcont
        RECT 6 20.5 8 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 7 25.5 dcont
        RECT 6 24.5 8 26.5 ;
      # VIA 2 21.5 dcont
        RECT 1 20.5 3 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 2 23.5 dcont
        RECT 1 22.5 3 24.5 ;
      # VIA 2 25.5 dcont
        RECT 1 24.5 3 26.5 ;
      # VIA 7 23.5 dcont
        RECT 6 22.5 8 24.5 ;
    END
END nr21
MACRO nr212
    CLASS core ;
    FOREIGN nr212 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 9.5 8.5 11.5 10.5 ;
        LAYER ML1 ;
        RECT 9.5 8.5 11.5 10.5 ;
        END
    END YB
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 8.5 6.0 10.5 ;
        LAYER ML1 ;
        RECT 4.0 8.5 6.0 10.5 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 11.5 9.0 13.5 ;
        LAYER ML1 ;
        RECT 7.0 11.5 9.0 13.5 ;
        END
    END B0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 1.5 24.5 1.5 18.0 7.5 18.0 7.5 24.5 ;
        WIDTH 2 ;
        PATH 4.5 21.5 4.5 28.5 ;
        
        
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 6.5 7.0 6.5 7.0 3.5 ;
        WIDTH 2 ;
        PATH 9.5 1.0 9.5 3.5 ;
        WIDTH 1.4 ;
        PATH 10.5 22.3 10.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 10.5 21.5 dcont
        RECT 9.5 20.5 11.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 10.5 25.5 dcont
        RECT 9.5 24.5 11.5 26.5 ;
      # VIA 6.5 3.5 dcont
        RECT 5.5 2.5 7.5 4.5 ;
      # VIA 9.5 3.5 dcont
        RECT 8.5 2.5 10.5 4.5 ;
      # VIA 10.5 23.5 dcont
        RECT 9.5 22.5 11.5 24.5 ;
    END
END nr212
MACRO nr222
    CLASS core ;
    FOREIGN nr222 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 12.5 8.0 14.5 10.0 ;
        LAYER ML1 ;
        RECT 12.5 8.0 14.5 10.0 ;
        END
    END YB
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.0 3.0 16.0 ;
        LAYER ML1 ;
        RECT 1.0 14.0 3.0 16.0 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 8.5 6.0 10.5 ;
        LAYER ML1 ;
        RECT 4.0 8.5 6.0 10.5 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 11.5 9.0 13.5 ;
        LAYER ML1 ;
        RECT 7.0 11.5 9.0 13.5 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 14.0 12.0 16.0 ;
        LAYER ML1 ;
        RECT 10.0 14.0 12.0 16.0 ;
        END
    END B0
    OBS
        LAYER ML1 ;
        
        WIDTH 2 ;
        PATH 11.5 1.0 11.5 3.5 ;
        WIDTH 1.4 ;
        PATH 10.5 20.0 10.5 24.0 ;
        WIDTH 1 ;
        PATH 10.5 20.5 10.5 17.5 13.5 17.5 13.5 6.5 7.0 6.5 7.0 3.5 ;
        WIDTH 1 ;
        PATH 1.5 24.0 1.5 17.5 7.5 17.5 7.5 26.5 13.5 26.5 13.5 20.0 ;
        
        
        WIDTH 2 ;
        PATH 4.5 20.0 4.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 1.5 20.8 1.5 24.0 ;
        
        LAYER ML1 ;
      # VIA 10.5 24 dcont
        RECT 9.5 23 11.5 25 ;
      # VIA 10.5 20 dcont
        RECT 9.5 19 11.5 21 ;
      # VIA 6.5 3.5 dcont
        RECT 5.5 2.5 7.5 4.5 ;
      # VIA 11.5 3.5 dcont
        RECT 10.5 2.5 12.5 4.5 ;
      # VIA 13.5 24 dcont
        RECT 12.5 23 14.5 25 ;
      # VIA 1.5 24 dcont
        RECT 0.5 23 2.5 25 ;
      # VIA 7.5 20 dcont
        RECT 6.5 19 8.5 21 ;
      # VIA 1.5 20 dcont
        RECT 0.5 19 2.5 21 ;
      # VIA 7.5 22 dcont
        RECT 6.5 21 8.5 23 ;
      # VIA 13.5 22 dcont
        RECT 12.5 21 14.5 23 ;
      # VIA 4.5 22 dcont
        RECT 3.5 21 5.5 23 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 13.5 20 dcont
        RECT 12.5 19 14.5 21 ;
      # VIA 10.5 22 dcont
        RECT 9.5 21 11.5 23 ;
      # VIA 7.5 24 dcont
        RECT 6.5 23 8.5 25 ;
      # VIA 4.5 20 dcont
        RECT 3.5 19 5.5 21 ;
      # VIA 1.5 22 dcont
        RECT 0.5 21 2.5 23 ;
      # VIA 4.5 24 dcont
        RECT 3.5 23 5.5 25 ;
    END
END nr222
MACRO nr31
    CLASS core ;
    FOREIGN nr31 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 8.0 12.0 10.0 ;
        LAYER ML1 ;
        RECT 10.0 8.0 12.0 10.0 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 12.0 9.0 14.0 ;
        LAYER ML1 ;
        RECT 7.0 12.0 9.0 14.0 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 9.5 20.5 9.5 18.0 10.5 18.0 10.5 3.6 ;
        WIDTH 1.4 ;
        PATH 9.5 22.3 9.5 25.5 ;
        WIDTH 1 ;
        PATH 5.0 3.5 5.0 6.5 10.5 6.5 ;
        WIDTH 2 ;
        PATH 7.5 1.0 7.5 3.8 ;
        
        
        WIDTH 2 ;
        PATH 2.5 21.5 2.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        
        LAYER ML1 ;
      # VIA 2.5 25.5 dcont
        RECT 1.5 24.5 3.5 26.5 ;
      # VIA 9.5 25.5 dcont
        RECT 8.5 24.5 10.5 26.5 ;
      # VIA 2.5 23.5 dcont
        RECT 1.5 22.5 3.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 9.5 21.5 dcont
        RECT 8.5 20.5 10.5 22.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 9.5 23.5 dcont
        RECT 8.5 22.5 10.5 24.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 2.5 21.5 dcont
        RECT 1.5 20.5 3.5 22.5 ;
    END
END nr31
MACRO or21
    CLASS core ;
    FOREIGN or21 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 12.5 BY 29.0 ;
    PIN Y
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.0 8.0 12.0 10.0 ;
        LAYER ML1 ;
        RECT 10.0 8.0 12.0 10.0 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 13.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 8.5 3.0 10.5 ;
        LAYER ML1 ;
        RECT 1.0 8.5 3.0 10.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 13.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 1.4 ;
        PATH 2.0 22.3 2.0 25.5 ;
        WIDTH 1 ;
        PATH 5.0 3.5 5.0 6.0 7.5 6.0 7.5 16.5 2.0 16.5 2.0 20.5 ;
        
        
        WIDTH 2 ;
        PATH 7.0 21.5 7.0 28.5 ;
        WIDTH 2 ;
        PATH 7.5 1.0 7.5 3.5 ;
        WIDTH 1.4 ;
        PATH 10.0 22.3 10.0 25.5 ;
        WIDTH 1 ;
        PATH 10.5 3.5 10.5 18.0 10.0 18.0 10.0 20.5 ;
        
        
        LAYER ML1 ;
      # VIA 7 23.5 dcont
        RECT 6 22.5 8 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7 21.5 dcont
        RECT 6 20.5 8 22.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 8 12.5 pcont
        RECT 7 11.5 9 13.5 ;
      # VIA 2 21.5 dcont
        RECT 1 20.5 3 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 10 23.5 dcont
        RECT 9 22.5 11 24.5 ;
      # VIA 2 23.5 dcont
        RECT 1 22.5 3 24.5 ;
      # VIA 10 21.5 dcont
        RECT 9 20.5 11 22.5 ;
      # VIA 2 25.5 dcont
        RECT 1 24.5 3 26.5 ;
      # VIA 7 25.5 dcont
        RECT 6 24.5 8 26.5 ;
      # VIA 10 25.5 dcont
        RECT 9 24.5 11 26.5 ;
    END
END or21
MACRO or31
    CLASS core ;
    FOREIGN or31 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 15.5 BY 29.0 ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 16.0 30.0 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.0 11.5 6.0 13.5 ;
        LAYER ML1 ;
        RECT 4.0 11.5 6.0 13.5 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.0 9.0 15.0 11.0 ;
        LAYER ML1 ;
        RECT 13.0 9.0 15.0 11.0 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.0 12.0 9.0 14.0 ;
        LAYER ML1 ;
        RECT 7.0 12.0 9.0 14.0 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 16.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 13.5 3.9 13.5 16.5 12.5 16.5 12.5 20.5 ;
        WIDTH 1.4 ;
        PATH 12.5 22.3 12.5 25.5 ;
        WIDTH 2 ;
        PATH 10.5 1.0 10.5 3.5 ;
        WIDTH 2 ;
        PATH 9.5 21.5 9.5 28.5 ;
        WIDTH 1 ;
        PATH 7.5 3.9 7.5 8.0 ;
        
        
        WIDTH 1 ;
        PATH 3.0 20.5 3.0 18.0 10.5 18.0 10.5 8.0 2.0 8.0 2.0 3.8 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.5 ;
        WIDTH 1.4 ;
        PATH 2.5 22.3 2.5 25.5 ;
        
        LAYER ML1 ;
      # VIA 9.5 25.5 dcont
        RECT 8.5 24.5 10.5 26.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 9.5 21.5 dcont
        RECT 8.5 20.5 10.5 22.5 ;
      # VIA 12.5 21.5 dcont
        RECT 11.5 20.5 13.5 22.5 ;
      # VIA 2.5 21.5 dcont
        RECT 1.5 20.5 3.5 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 10.5 3.5 dcont
        RECT 9.5 2.5 11.5 4.5 ;
      # VIA 2.5 25.5 dcont
        RECT 1.5 24.5 3.5 26.5 ;
      # VIA 12.5 25.5 dcont
        RECT 11.5 24.5 13.5 26.5 ;
      # VIA 2.5 23.5 dcont
        RECT 1.5 22.5 3.5 24.5 ;
      # VIA 11 13 pcont
        RECT 10 12 12 14 ;
      # VIA 9.5 23.5 dcont
        RECT 8.5 22.5 10.5 24.5 ;
      # VIA 12.5 23.5 dcont
        RECT 11.5 22.5 13.5 24.5 ;
      # VIA 13.5 3.5 dcont
        RECT 12.5 2.5 14.5 4.5 ;
    END
END or31
MACRO rff1
    CLASS core ;
    FOREIGN rff1 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 56.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN R
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 43.0 10.5 45.0 12.5 ;
        LAYER ML1 ;
        RECT 43.0 10.5 45.0 12.5 ;
        END
    END R
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 53.5 10.5 55.5 12.5 ;
        LAYER ML1 ;
        RECT 53.5 10.5 55.5 12.5 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 56.5 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 56.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 1.5 26.0 1.5 3.6 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 5.4 13.0 1.5 13.0 ;
        WIDTH 1 ;
        PATH 5.9 19.0 1.8 19.0 ;
        WIDTH 1 ;
        PATH 5.9 6.5 1.5 6.5 ;
        WIDTH 2 ;
        PATH 4.5 22.6 4.5 28.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.8 ;
        WIDTH 1 ;
        PATH 8.0 3.6 8.0 9.5 7.5 9.5 7.5 16.0 8.0 16.0 8.0 26.0 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 1 ;
        PATH 14.9 6.5 8.0 6.5 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 16.0 22.6 16.0 19.0 22.3 19.0 ;
        WIDTH 1 ;
        PATH 16.3 3.8 16.3 4.0 17.5 4.0 17.5 10.0 22.4 10.0 ;
        WIDTH 1 ;
        PATH 7.5 16.0 32.0 16.0 ;
        WIDTH 2 ;
        PATH 21.0 22.6 21.0 28.5 ;
        WIDTH 2 ;
        PATH 21.0 1.0 21.0 3.8 ;
        WIDTH 1 ;
        PATH 36.0 13.0 10.3 13.0 ;
        WIDTH 1 ;
        PATH 28.3 6.5 19.9 6.5 ;
        WIDTH 1 ;
        PATH 24.0 3.8 24.0 6.5 ;
        WIDTH 1.4 ;
        PATH 26.0 22.3 26.0 25.5 ;
        WIDTH 2 ;
        PATH 27.0 1.0 27.0 3.8 ;
        WIDTH 1 ;
        PATH 26.0 22.6 26.0 19.0 28.3 19.0 ;
        
        
        WIDTH 2 ;
        PATH 29.5 22.6 29.5 28.5 ;
        WIDTH 1 ;
        PATH 25.5 10.0 44.5 10.0 ;
        WIDTH 1.4 ;
        PATH 34.5 22.3 34.5 25.5 ;
        WIDTH 1 ;
        PATH 32.5 3.8 32.5 6.0 37.8 6.0 ;
        WIDTH 2 ;
        PATH 37.0 1.0 37.0 3.8 ;
        WIDTH 1 ;
        PATH 34.5 22.6 34.5 19.0 41.0 19.0 ;
        WIDTH 2 ;
        PATH 39.5 22.6 39.5 28.5 ;
        WIDTH 1 ;
        PATH 38.5 14.0 44.9 14.0 ;
        WIDTH 2 ;
        PATH 43.0 1.0 43.0 3.8 ;
        WIDTH 1.4 ;
        PATH 44.5 22.3 44.5 25.5 ;
        WIDTH 1 ;
        PATH 40.5 3.8 40.5 6.0 46.5 6.0 46.5 8.5 48.5 8.5 48.5 14.0 44.5 14.0 44.5 21.5 ;
        WIDTH 1 ;
        PATH 49.3 16.5 44.5 16.5 ;
        WIDTH 1.4 ;
        PATH 48.0 22.3 48.0 25.5 ;
        WIDTH 1 ;
        PATH 48.0 26.0 48.0 19.0 52.0 19.0 52.0 6.0 48.5 6.0 48.5 3.6 ;
        WIDTH 2 ;
        PATH 51.0 1.0 51.0 3.8 ;
        WIDTH 2 ;
        PATH 51.0 22.6 51.0 28.5 ;
        WIDTH 1.4 ;
        PATH 54.0 22.3 54.0 25.5 ;
        WIDTH 1 ;
        PATH 54.5 3.3 54.5 26.0 ;
        
        LAYER ML1 ;
      # VIA 40.5 18.5 pcont
        RECT 39.5 17.5 41.5 19.5 ;
      # VIA 40 3.5 dcont
        RECT 39 2.5 41 4.5 ;
      # VIA 26 25.5 dcont
        RECT 25 24.5 27 26.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 43 3.5 dcont
        RECT 42 2.5 44 4.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 39.5 25.5 dcont
        RECT 38.5 24.5 40.5 26.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 38.5 14 pcont
        RECT 37.5 13 39.5 15 ;
      # VIA 26 23.5 dcont
        RECT 25 22.5 27 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 48 3.5 dcont
        RECT 47 2.5 49 4.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 49 16.5 pcont
        RECT 48 15.5 50 17.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 54 21.5 dcont
        RECT 53 20.5 55 22.5 ;
      # VIA 39.5 21.5 dcont
        RECT 38.5 20.5 40.5 22.5 ;
      # VIA 29.5 25.5 dcont
        RECT 28.5 24.5 30.5 26.5 ;
      # VIA 54 3.5 dcont
        RECT 53 2.5 55 4.5 ;
      # VIA 48 25.5 dcont
        RECT 47 24.5 49 26.5 ;
      # VIA 34.5 23.5 dcont
        RECT 33.5 22.5 35.5 24.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 34.5 25.5 dcont
        RECT 33.5 24.5 35.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 44.5 21.5 dcont
        RECT 43.5 20.5 45.5 22.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 38 6.5 pcont
        RECT 37 5.5 39 7.5 ;
      # VIA 28 18.5 pcont
        RECT 27 17.5 29 19.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 20 6.5 pcont
        RECT 19 5.5 21 7.5 ;
      # VIA 44.5 23.5 dcont
        RECT 43.5 22.5 45.5 24.5 ;
      # VIA 48 21.5 dcont
        RECT 47 20.5 49 22.5 ;
      # VIA 52 18.5 pcont
        RECT 51 17.5 53 19.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 54 23.5 dcont
        RECT 53 22.5 55 24.5 ;
      # VIA 27 3.5 dcont
        RECT 26 2.5 28 4.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 54 25.5 dcont
        RECT 53 24.5 55 26.5 ;
      # VIA 44.5 25.5 dcont
        RECT 43.5 24.5 45.5 26.5 ;
      # VIA 26 21.5 dcont
        RECT 25 20.5 27 22.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 34.5 21.5 dcont
        RECT 33.5 20.5 35.5 22.5 ;
      # VIA 32 16.5 pcont
        RECT 31 15.5 33 17.5 ;
      # VIA 39.5 23.5 dcont
        RECT 38.5 22.5 40.5 24.5 ;
      # VIA 49 9 pcont
        RECT 48 8 50 10 ;
      # VIA 52 6.5 pcont
        RECT 51 5.5 53 7.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 30 13 pcont
        RECT 29 12 31 14 ;
      # VIA 35.5 14 pcont
        RECT 34.5 13 36.5 15 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 24 3.5 dcont
        RECT 23 2.5 25 4.5 ;
      # VIA 32 3.5 dcont
        RECT 31 2.5 33 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 37 3.5 dcont
        RECT 36 2.5 38 4.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 25 10 pcont
        RECT 24 9 26 11 ;
      # VIA 48 23.5 dcont
        RECT 47 22.5 49 24.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 29.5 21.5 dcont
        RECT 28.5 20.5 30.5 22.5 ;
      # VIA 29.5 23.5 dcont
        RECT 28.5 22.5 30.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 28 6.5 pcont
        RECT 27 5.5 29 7.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 15 13 pcont
        RECT 14 12 16 14 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
    END
END rff1
MACRO rff1_r
    CLASS core ;
    FOREIGN rff1_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 62.5 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN R
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.5 51.5 12.5 ;
        LAYER ML1 ;
        RECT 49.5 10.5 51.5 12.5 ;
        END
    END R
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 60.0 10.5 62.0 12.5 ;
        LAYER ML1 ;
        RECT 60.0 10.5 62.0 12.5 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 63.0 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 63.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 61.0 3.3 61.0 26.0 ;
        WIDTH 1.4 ;
        PATH 60.5 22.3 60.5 25.5 ;
        WIDTH 2 ;
        PATH 57.5 22.6 57.5 28.5 ;
        WIDTH 2 ;
        PATH 57.5 1.0 57.5 3.8 ;
        WIDTH 1 ;
        PATH 54.5 26.0 54.5 19.0 58.5 19.0 58.5 6.0 55.0 6.0 55.0 3.6 ;
        WIDTH 1.4 ;
        PATH 54.5 22.3 54.5 25.5 ;
        WIDTH 1 ;
        PATH 55.8 16.5 51.0 16.5 ;
        WIDTH 1 ;
        PATH 47.0 3.8 47.0 6.0 53.0 6.0 53.0 8.5 55.0 8.5 55.0 14.0 51.0 14.0 51.0 21.5 ;
        WIDTH 1.4 ;
        PATH 51.0 22.3 51.0 25.5 ;
        WIDTH 2 ;
        PATH 49.5 1.0 49.5 3.8 ;
        WIDTH 1 ;
        PATH 45.0 14.0 51.4 14.0 ;
        WIDTH 2 ;
        PATH 46.0 22.6 46.0 28.5 ;
        WIDTH 1 ;
        PATH 41.0 22.6 41.0 19.0 47.5 19.0 ;
        WIDTH 2 ;
        PATH 43.5 1.0 43.5 3.8 ;
        WIDTH 1 ;
        PATH 39.0 3.8 39.0 6.0 44.3 6.0 ;
        WIDTH 1.4 ;
        PATH 41.0 22.3 41.0 25.5 ;
        WIDTH 1 ;
        PATH 32.0 10.0 51.0 10.0 ;
        WIDTH 2 ;
        PATH 36.0 22.6 36.0 28.5 ;
        
        
        WIDTH 1 ;
        PATH 32.5 22.6 32.5 19.0 34.8 19.0 ;
        WIDTH 2 ;
        PATH 33.5 1.0 33.5 3.8 ;
        WIDTH 1.4 ;
        PATH 32.5 22.3 32.5 25.5 ;
        WIDTH 1 ;
        PATH 30.5 3.8 30.5 6.5 ;
        WIDTH 1 ;
        PATH 34.8 6.5 26.4 6.5 ;
        WIDTH 1 ;
        PATH 42.5 13.0 16.8 13.0 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.8 ;
        WIDTH 2 ;
        PATH 27.5 22.6 27.5 28.5 ;
        WIDTH 1 ;
        PATH 14.0 16.0 38.5 16.0 ;
        WIDTH 1 ;
        PATH 22.8 3.8 22.8 4.0 24.0 4.0 24.0 10.0 28.9 10.0 ;
        WIDTH 1 ;
        PATH 22.5 22.6 22.5 19.0 28.8 19.0 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 21.4 6.5 14.5 6.5 ;
        WIDTH 2 ;
        PATH 17.5 22.6 17.5 28.5 ;
        WIDTH 2 ;
        PATH 17.5 1.0 17.5 3.8 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 16.0 14.5 16.0 14.5 26.0 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 1 ;
        PATH 12.4 6.5 8.0 6.5 ;
        WIDTH 1 ;
        PATH 12.4 19.0 8.3 19.0 ;
        WIDTH 1 ;
        PATH 11.9 13.0 8.0 13.0 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 8.0 26.0 8.0 3.6 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        
        LAYER ML1 ;
      # VIA 5.5 13 pcont
        RECT 4.5 12 6.5 14 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 34.5 6.5 pcont
        RECT 33.5 5.5 35.5 7.5 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 36 23.5 dcont
        RECT 35 22.5 37 24.5 ;
      # VIA 36 21.5 dcont
        RECT 35 20.5 37 22.5 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 54.5 23.5 dcont
        RECT 53.5 22.5 55.5 24.5 ;
      # VIA 31.5 10 pcont
        RECT 30.5 9 32.5 11 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 43.5 3.5 dcont
        RECT 42.5 2.5 44.5 4.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 38.5 3.5 dcont
        RECT 37.5 2.5 39.5 4.5 ;
      # VIA 30.5 3.5 dcont
        RECT 29.5 2.5 31.5 4.5 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 42 14 pcont
        RECT 41 13 43 15 ;
      # VIA 36.5 13 pcont
        RECT 35.5 12 37.5 14 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 55.5 9 pcont
        RECT 54.5 8 56.5 10 ;
      # VIA 58.5 6.5 pcont
        RECT 57.5 5.5 59.5 7.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 46 23.5 dcont
        RECT 45 22.5 47 24.5 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 38.5 16.5 pcont
        RECT 37.5 15.5 39.5 17.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 41 21.5 dcont
        RECT 40 20.5 42 22.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 32.5 21.5 dcont
        RECT 31.5 20.5 33.5 22.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 60.5 25.5 dcont
        RECT 59.5 24.5 61.5 26.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 57.5 23.5 dcont
        RECT 56.5 22.5 58.5 24.5 ;
      # VIA 33.5 3.5 dcont
        RECT 32.5 2.5 34.5 4.5 ;
      # VIA 60.5 23.5 dcont
        RECT 59.5 22.5 61.5 24.5 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 58.5 18.5 pcont
        RECT 57.5 17.5 59.5 19.5 ;
      # VIA 54.5 21.5 dcont
        RECT 53.5 20.5 55.5 22.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 34.5 18.5 pcont
        RECT 33.5 17.5 35.5 19.5 ;
      # VIA 44.5 6.5 pcont
        RECT 43.5 5.5 45.5 7.5 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 41 25.5 dcont
        RECT 40 24.5 42 26.5 ;
      # VIA 57.5 25.5 dcont
        RECT 56.5 24.5 58.5 26.5 ;
      # VIA 41 23.5 dcont
        RECT 40 22.5 42 24.5 ;
      # VIA 54.5 25.5 dcont
        RECT 53.5 24.5 55.5 26.5 ;
      # VIA 60.5 3.5 dcont
        RECT 59.5 2.5 61.5 4.5 ;
      # VIA 36 25.5 dcont
        RECT 35 24.5 37 26.5 ;
      # VIA 46 21.5 dcont
        RECT 45 20.5 47 22.5 ;
      # VIA 60.5 21.5 dcont
        RECT 59.5 20.5 61.5 22.5 ;
      # VIA 28.5 10 pcont
        RECT 27.5 9 29.5 11 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 55.5 16.5 pcont
        RECT 54.5 15.5 56.5 17.5 ;
      # VIA 57.5 21.5 dcont
        RECT 56.5 20.5 58.5 22.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 54.5 3.5 dcont
        RECT 53.5 2.5 55.5 4.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 21.5 13 pcont
        RECT 20.5 12 22.5 14 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 32.5 23.5 dcont
        RECT 31.5 22.5 33.5 24.5 ;
      # VIA 45 14 pcont
        RECT 44 13 46 15 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 46 25.5 dcont
        RECT 45 24.5 47 26.5 ;
      # VIA 57.5 3.5 dcont
        RECT 56.5 2.5 58.5 4.5 ;
      # VIA 49.5 3.5 dcont
        RECT 48.5 2.5 50.5 4.5 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 32.5 25.5 dcont
        RECT 31.5 24.5 33.5 26.5 ;
      # VIA 46.5 3.5 dcont
        RECT 45.5 2.5 47.5 4.5 ;
      # VIA 47 18.5 pcont
        RECT 46 17.5 48 19.5 ;
    END
END rff1_r
MACRO rff1m2
    CLASS core ;
    FOREIGN rff1m2 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 56.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCk ;
        PORT
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN R
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 43.0 10.5 45.0 12.5 ;
        LAYER ML2 ;
        RECT 43.0 10.5 45.0 12.5 ;
        END
    END R
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 53.5 10.5 55.5 12.5 ;
        LAYER ML2 ;
        RECT 53.5 10.5 55.5 12.5 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 56.5 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 56.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 1.5 26.0 1.5 3.6 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 5.4 13.0 1.5 13.0 ;
        WIDTH 1 ;
        PATH 5.6 18.5 1.5 18.5 ;
        WIDTH 1 ;
        PATH 5.9 6.5 1.5 6.5 ;
        WIDTH 2 ;
        PATH 4.5 22.6 4.5 28.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.8 ;
        WIDTH 1 ;
        PATH 8.0 3.6 8.0 9.5 7.5 9.5 7.5 16.0 8.0 16.0 8.0 26.0 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 1 ;
        PATH 14.8 6.5 8.3 6.5 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 16.0 22.6 16.0 19.0 22.3 19.0 ;
        WIDTH 1 ;
        PATH 16.3 3.8 16.3 4.0 17.5 4.0 17.5 10.0 22.4 10.0 ;
        WIDTH 1 ;
        PATH 7.5 16.0 33.3 16.0 ;
        WIDTH 2 ;
        PATH 21.0 22.6 21.0 28.5 ;
        WIDTH 2 ;
        PATH 21.0 1.0 21.0 3.8 ;
        WIDTH 1 ;
        PATH 35.8 13.0 10.3 13.0 ;
        WIDTH 1 ;
        PATH 28.3 6.5 19.9 6.5 ;
        WIDTH 1 ;
        PATH 24.0 3.8 24.0 6.5 ;
        WIDTH 1.4 ;
        PATH 26.0 22.3 26.0 25.5 ;
        WIDTH 2 ;
        PATH 27.0 1.0 27.0 3.8 ;
        WIDTH 1 ;
        PATH 26.0 22.6 26.0 19.0 28.3 19.0 ;
        
        
        WIDTH 2 ;
        PATH 29.5 22.6 29.5 28.5 ;
        WIDTH 1 ;
        PATH 25.4 10.0 44.5 10.0 ;
        WIDTH 1.4 ;
        PATH 34.5 22.3 34.5 25.5 ;
        WIDTH 1 ;
        PATH 32.5 3.8 32.5 6.5 37.8 6.5 ;
        WIDTH 2 ;
        PATH 37.0 1.0 37.0 3.8 ;
        WIDTH 1 ;
        PATH 34.5 22.6 34.5 19.0 41.0 19.0 ;
        WIDTH 2 ;
        PATH 39.5 22.6 39.5 28.5 ;
        WIDTH 1 ;
        PATH 38.5 14.0 44.9 14.0 ;
        WIDTH 2 ;
        PATH 43.0 1.0 43.0 3.8 ;
        WIDTH 1.4 ;
        PATH 44.5 22.3 44.5 25.5 ;
        WIDTH 1 ;
        PATH 40.5 3.8 40.5 6.0 46.5 6.0 46.5 8.5 48.5 8.5 48.5 14.0 45.0 14.0 45.0 21.5 ;
        WIDTH 1 ;
        PATH 49.3 17.0 45.0 17.0 ;
        WIDTH 1.4 ;
        PATH 48.0 22.3 48.0 25.5 ;
        WIDTH 1 ;
        PATH 48.5 26.0 48.5 19.0 52.0 19.0 52.0 6.0 48.5 6.0 48.5 3.6 ;
        WIDTH 2 ;
        PATH 51.0 1.0 51.0 3.8 ;
        WIDTH 2 ;
        PATH 51.0 22.6 51.0 28.5 ;
        RECT 53 2.5 55 4.5 ;
        WIDTH 1.4 ;
        PATH 54.0 22.3 54.0 25.5 ;
        WIDTH 1 ;
        PATH 54.5 3.3 54.5 26.0 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 22.0 10.0 22.0 18.7 ;
        WIDTH 1 ;
        PATH 28.0 18.6 28.0 6.8 ;
        WIDTH 1 ;
        PATH 40.0 18.6 40.0 16.0 38.5 16.0 38.5 6.8 ;
        LAYER ML1 ;
      # VIA 40.5 18.5 pcont
        RECT 39.5 17.5 41.5 19.5 ;
      # VIA 40 3.5 dcont
        RECT 39 2.5 41 4.5 ;
      # VIA 26 25.5 dcont
        RECT 25 24.5 27 26.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 43 3.5 dcont
        RECT 42 2.5 44 4.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 39.5 25.5 dcont
        RECT 38.5 24.5 40.5 26.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 38.5 14 pcont
        RECT 37.5 13 39.5 15 ;
      # VIA 26 23.5 dcont
        RECT 25 22.5 27 24.5 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML2 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML1 ;
      # VIA 48 3.5 dcont
        RECT 47 2.5 49 4.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 49 16.5 pcont
        RECT 48 15.5 50 17.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 54 21.5 dcont
        RECT 53 20.5 55 22.5 ;
      # VIA 39.5 21.5 dcont
        RECT 38.5 20.5 40.5 22.5 ;
      # VIA 29.5 25.5 dcont
        RECT 28.5 24.5 30.5 26.5 ;
      # VIA 54 3.5 dcont
        RECT 53 2.5 55 4.5 ;
      # VIA 48 25.5 dcont
        RECT 47 24.5 49 26.5 ;
      # VIA 34.5 23.5 dcont
        RECT 33.5 22.5 35.5 24.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 34.5 25.5 dcont
        RECT 33.5 24.5 35.5 26.5 ;
      # VIA 28 7 dcont
        RECT 27 6 29 8 ;
        LAYER ML2 ;
      # VIA 28 7 dcont
        RECT 27 6 29 8 ;
        LAYER ML1 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 44.5 21.5 dcont
        RECT 43.5 20.5 45.5 22.5 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
      # VIA 38 7 pcont
        RECT 37 6 39 8 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 15 13 pcont
        RECT 14 12 16 14 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 20 7 pcont
        RECT 19 6 21 8 ;
      # VIA 44.5 23.5 dcont
        RECT 43.5 22.5 45.5 24.5 ;
      # VIA 48 21.5 dcont
        RECT 47 20.5 49 22.5 ;
      # VIA 52 18.5 pcont
        RECT 51 17.5 53 19.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML2 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML1 ;
      # VIA 54 23.5 dcont
        RECT 53 22.5 55 24.5 ;
      # VIA 27 3.5 dcont
        RECT 26 2.5 28 4.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 54 25.5 dcont
        RECT 53 24.5 55 26.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 44.5 25.5 dcont
        RECT 43.5 24.5 45.5 26.5 ;
      # VIA 26 21.5 dcont
        RECT 25 20.5 27 22.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 34.5 21.5 dcont
        RECT 33.5 20.5 35.5 22.5 ;
      # VIA 33 16.5 pcont
        RECT 32 15.5 34 17.5 ;
      # VIA 39.5 23.5 dcont
        RECT 38.5 22.5 40.5 24.5 ;
      # VIA 38 7 dcont
        RECT 37 6 39 8 ;
        LAYER ML2 ;
      # VIA 38 7 dcont
        RECT 37 6 39 8 ;
        LAYER ML1 ;
      # VIA 52 6.5 pcont
        RECT 51 5.5 53 7.5 ;
      # VIA 49 9 pcont
        RECT 48 8 50 10 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 30 13 pcont
        RECT 29 12 31 14 ;
      # VIA 40.5 18.5 dcont
        RECT 39.5 17.5 41.5 19.5 ;
        LAYER ML2 ;
      # VIA 40.5 18.5 dcont
        RECT 39.5 17.5 41.5 19.5 ;
        LAYER ML1 ;
      # VIA 35.5 13.5 pcont
        RECT 34.5 12.5 36.5 14.5 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML2 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML1 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 24 3.5 dcont
        RECT 23 2.5 25 4.5 ;
      # VIA 32 3.5 dcont
        RECT 31 2.5 33 4.5 ;
      # VIA 37 3.5 dcont
        RECT 36 2.5 38 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 25.5 10 pcont
        RECT 24.5 9 26.5 11 ;
      # VIA 48 23.5 dcont
        RECT 47 22.5 49 24.5 ;
      # VIA 29.5 21.5 dcont
        RECT 28.5 20.5 30.5 22.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 29.5 23.5 dcont
        RECT 28.5 22.5 30.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 28 7 pcont
        RECT 27 6 29 8 ;
    END
END rff1m2
MACRO rff1m2_r
    CLASS core ;
    FOREIGN rff1m2_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 62.5 BY 29.0 ;
    PIN R
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.5 51.5 12.5 ;
        LAYER ML1 ;
        RECT 49.5 10.5 51.5 12.5 ;
        END
    END R
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 63.0 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 60.0 10.5 62.0 12.5 ;
        LAYER ML1 ;
        RECT 60.0 10.5 62.0 12.5 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 63.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 8.0 26.0 8.0 3.6 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 11.9 13.0 8.0 13.0 ;
        WIDTH 1 ;
        PATH 12.1 18.5 8.0 18.5 ;
        WIDTH 1 ;
        PATH 12.4 6.5 8.0 6.5 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 16.0 14.5 16.0 14.5 26.0 ;
        WIDTH 2 ;
        PATH 17.5 1.0 17.5 3.8 ;
        WIDTH 2 ;
        PATH 17.5 22.6 17.5 28.5 ;
        WIDTH 1 ;
        PATH 21.3 6.5 14.8 6.5 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 22.5 22.6 22.5 19.0 28.8 19.0 ;
        WIDTH 1 ;
        PATH 22.8 3.8 22.8 4.0 24.0 4.0 24.0 10.0 28.9 10.0 ;
        WIDTH 1 ;
        PATH 14.0 16.0 39.8 16.0 ;
        WIDTH 2 ;
        PATH 27.5 22.6 27.5 28.5 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.8 ;
        WIDTH 1 ;
        PATH 42.3 13.0 16.8 13.0 ;
        WIDTH 1 ;
        PATH 34.8 6.5 26.4 6.5 ;
        WIDTH 1 ;
        PATH 30.5 3.8 30.5 6.5 ;
        WIDTH 1.4 ;
        PATH 32.5 22.3 32.5 25.5 ;
        WIDTH 2 ;
        PATH 33.5 1.0 33.5 3.8 ;
        WIDTH 1 ;
        PATH 32.5 22.6 32.5 19.0 34.8 19.0 ;
        
        
        WIDTH 2 ;
        PATH 36.0 22.6 36.0 28.5 ;
        WIDTH 1 ;
        PATH 31.9 10.0 51.0 10.0 ;
        WIDTH 1.4 ;
        PATH 41.0 22.3 41.0 25.5 ;
        WIDTH 1 ;
        PATH 39.0 3.8 39.0 6.5 44.3 6.5 ;
        WIDTH 2 ;
        PATH 43.5 1.0 43.5 3.8 ;
        WIDTH 1 ;
        PATH 41.0 22.6 41.0 19.0 47.5 19.0 ;
        WIDTH 2 ;
        PATH 46.0 22.6 46.0 28.5 ;
        WIDTH 1 ;
        PATH 45.0 14.0 51.4 14.0 ;
        WIDTH 2 ;
        PATH 49.5 1.0 49.5 3.8 ;
        WIDTH 1.4 ;
        PATH 51.0 22.3 51.0 25.5 ;
        WIDTH 1 ;
        PATH 47.0 3.8 47.0 6.0 53.0 6.0 53.0 8.5 55.0 8.5 55.0 14.0 51.5 14.0 51.5 21.5 ;
        WIDTH 1 ;
        PATH 55.8 17.0 51.5 17.0 ;
        WIDTH 1.4 ;
        PATH 54.5 22.3 54.5 25.5 ;
        WIDTH 1 ;
        PATH 55.0 26.0 55.0 19.0 58.5 19.0 58.5 6.0 55.0 6.0 55.0 3.6 ;
        WIDTH 2 ;
        PATH 57.5 1.0 57.5 3.8 ;
        WIDTH 2 ;
        PATH 57.5 22.6 57.5 28.5 ;
        RECT 59.5 2.5 61.5 4.5 ;
        WIDTH 1.4 ;
        PATH 60.5 22.3 60.5 25.5 ;
        WIDTH 1 ;
        PATH 61.0 3.3 61.0 26.0 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        
        
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 28.5 10.0 28.5 18.7 ;
        WIDTH 1 ;
        PATH 34.5 18.6 34.5 6.8 ;
        WIDTH 1 ;
        PATH 46.5 18.6 46.5 16.0 45.0 16.0 45.0 6.8 ;
        LAYER ML1 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 47 18.5 pcont
        RECT 46 17.5 48 19.5 ;
      # VIA 46.5 3.5 dcont
        RECT 45.5 2.5 47.5 4.5 ;
      # VIA 32.5 25.5 dcont
        RECT 31.5 24.5 33.5 26.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 49.5 3.5 dcont
        RECT 48.5 2.5 50.5 4.5 ;
      # VIA 57.5 3.5 dcont
        RECT 56.5 2.5 58.5 4.5 ;
      # VIA 46 25.5 dcont
        RECT 45 24.5 47 26.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 45 14 pcont
        RECT 44 13 46 15 ;
      # VIA 32.5 23.5 dcont
        RECT 31.5 22.5 33.5 24.5 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 35 18.5 dcont
        RECT 34 17.5 36 19.5 ;
        LAYER ML2 ;
      # VIA 35 18.5 dcont
        RECT 34 17.5 36 19.5 ;
        LAYER ML1 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 54.5 3.5 dcont
        RECT 53.5 2.5 55.5 4.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 57.5 21.5 dcont
        RECT 56.5 20.5 58.5 22.5 ;
      # VIA 55.5 16.5 pcont
        RECT 54.5 15.5 56.5 17.5 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 28.5 10 pcont
        RECT 27.5 9 29.5 11 ;
      # VIA 60.5 21.5 dcont
        RECT 59.5 20.5 61.5 22.5 ;
      # VIA 46 21.5 dcont
        RECT 45 20.5 47 22.5 ;
      # VIA 36 25.5 dcont
        RECT 35 24.5 37 26.5 ;
      # VIA 60.5 3.5 dcont
        RECT 59.5 2.5 61.5 4.5 ;
      # VIA 54.5 25.5 dcont
        RECT 53.5 24.5 55.5 26.5 ;
      # VIA 41 23.5 dcont
        RECT 40 22.5 42 24.5 ;
      # VIA 57.5 25.5 dcont
        RECT 56.5 24.5 58.5 26.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 41 25.5 dcont
        RECT 40 24.5 42 26.5 ;
      # VIA 34.5 7 dcont
        RECT 33.5 6 35.5 8 ;
        LAYER ML2 ;
      # VIA 34.5 7 dcont
        RECT 33.5 6 35.5 8 ;
        LAYER ML1 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 44.5 7 pcont
        RECT 43.5 6 45.5 8 ;
      # VIA 35 18.5 pcont
        RECT 34 17.5 36 19.5 ;
      # VIA 21.5 13 pcont
        RECT 20.5 12 22.5 14 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 26.5 7 pcont
        RECT 25.5 6 27.5 8 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 54.5 21.5 dcont
        RECT 53.5 20.5 55.5 22.5 ;
      # VIA 58.5 18.5 pcont
        RECT 57.5 17.5 59.5 19.5 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML2 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML1 ;
      # VIA 60.5 23.5 dcont
        RECT 59.5 22.5 61.5 24.5 ;
      # VIA 33.5 3.5 dcont
        RECT 32.5 2.5 34.5 4.5 ;
      # VIA 57.5 23.5 dcont
        RECT 56.5 22.5 58.5 24.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 60.5 25.5 dcont
        RECT 59.5 24.5 61.5 26.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 32.5 21.5 dcont
        RECT 31.5 20.5 33.5 22.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 41 21.5 dcont
        RECT 40 20.5 42 22.5 ;
      # VIA 39.5 16.5 pcont
        RECT 38.5 15.5 40.5 17.5 ;
      # VIA 46 23.5 dcont
        RECT 45 22.5 47 24.5 ;
      # VIA 44.5 7 dcont
        RECT 43.5 6 45.5 8 ;
        LAYER ML2 ;
      # VIA 44.5 7 dcont
        RECT 43.5 6 45.5 8 ;
        LAYER ML1 ;
      # VIA 58.5 6.5 pcont
        RECT 57.5 5.5 59.5 7.5 ;
      # VIA 55.5 9 pcont
        RECT 54.5 8 56.5 10 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 36.5 13 pcont
        RECT 35.5 12 37.5 14 ;
      # VIA 47 18.5 dcont
        RECT 46 17.5 48 19.5 ;
        LAYER ML2 ;
      # VIA 47 18.5 dcont
        RECT 46 17.5 48 19.5 ;
        LAYER ML1 ;
      # VIA 42 13.5 pcont
        RECT 41 12.5 43 14.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML2 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML1 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 30.5 3.5 dcont
        RECT 29.5 2.5 31.5 4.5 ;
      # VIA 38.5 3.5 dcont
        RECT 37.5 2.5 39.5 4.5 ;
      # VIA 43.5 3.5 dcont
        RECT 42.5 2.5 44.5 4.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 32 10 pcont
        RECT 31 9 33 11 ;
      # VIA 54.5 23.5 dcont
        RECT 53.5 22.5 55.5 24.5 ;
      # VIA 36 21.5 dcont
        RECT 35 20.5 37 22.5 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 36 23.5 dcont
        RECT 35 22.5 37 24.5 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 34.5 7 pcont
        RECT 33.5 6 35.5 8 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 5.5 13 pcont
        RECT 4.5 12 6.5 14 ;
    END
END rff1m2_r
MACRO sff1
    CLASS core ;
    FOREIGN sff1 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 56.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN S
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER ML2 ;
        RECT 43.0 10.0 45.0 12.0 ;
        LAYER ML1 ;
        RECT 43.0 10.0 45.0 12.0 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 53.5 10.5 55.5 12.5 ;
        LAYER ML1 ;
        RECT 53.5 10.5 55.5 12.5 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 56.5 30.0 ;
        END
    END VDD
    PIN VSS
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 56.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 24.5 19.0 24.5 21.5 ;
        WIDTH 1 ;
        PATH 31.8 15.5 7.8 15.5 ;
        WIDTH 0 ;
        PATH 44.0 10.8 44.0 9.3 25.3 9.3 ;
        WIDTH 0 ;
        PATH 44.0 10.8 44.0 9.3 25.3 9.3 ;
        WIDTH 1 ;
        PATH 1.5 26.0 1.5 3.6 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 5.4 13.0 1.5 13.0 ;
        WIDTH 1 ;
        PATH 5.8 6.0 1.5 6.0 ;
        WIDTH 1 ;
        PATH 5.6 18.5 1.5 18.5 ;
        WIDTH 2 ;
        PATH 4.5 22.6 4.5 28.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.8 ;
        RECT 6.9 20.9 8.1 26.1 ;
        WIDTH 1 ;
        PATH 8.0 3.6 8.0 9.5 7.5 9.5 7.5 15.5 8.0 15.5 8.0 26.0 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 1 ;
        PATH 14.8 6.5 8.3 6.5 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 16.0 22.3 16.0 19.0 22.0 19.0 ;
        WIDTH 1 ;
        PATH 16.0 3.8 16.0 4.0 17.5 4.0 17.5 9.5 22.1 9.5 ;
        WIDTH 2 ;
        PATH 21.0 22.6 21.0 28.5 ;
        WIDTH 2 ;
        PATH 21.0 1.0 21.0 3.8 ;
        WIDTH 1 ;
        PATH 35.4 12.5 10.3 12.5 ;
        WIDTH 1 ;
        PATH 27.3 6.0 20.3 6.0 ;
        WIDTH 1.4 ;
        PATH 24.0 21.5 24.0 25.5 ;
        WIDTH 1 ;
        PATH 24.5 19.0 28.5 19.0 28.5 18.0 ;
        WIDTH 1 ;
        PATH 26.5 3.6 26.5 5.5 ;
        WIDTH 2 ;
        PATH 27.0 23.8 27.0 28.5 ;
        
        
        WIDTH 2 ;
        PATH 29.5 1.0 29.5 3.8 ;
        WIDTH 1.4 ;
        PATH 33.5 22.3 33.5 25.5 ;
        WIDTH 1 ;
        PATH 34.0 22.3 34.0 19.0 39.5 19.0 ;
        WIDTH 2 ;
        PATH 38.5 22.6 38.5 28.5 ;
        WIDTH 1 ;
        PATH 35.0 3.8 35.0 6.0 40.3 6.0 ;
        WIDTH 2 ;
        PATH 39.5 1.0 39.5 3.8 ;
        WIDTH 2 ;
        PATH 44.5 22.6 44.5 28.5 ;
        WIDTH 1 ;
        PATH 45.0 3.8 45.0 8.0 49.5 8.0 49.5 17.0 42.3 17.0 ;
        WIDTH 1.4 ;
        PATH 48.0 22.3 48.0 25.5 ;
        WIDTH 1 ;
        PATH 48.5 26.0 48.5 19.0 52.0 19.0 52.0 6.0 48.5 6.0 48.5 3.6 ;
        WIDTH 2 ;
        PATH 51.0 1.0 51.0 3.8 ;
        WIDTH 2 ;
        PATH 51.0 22.6 51.0 28.5 ;
        WIDTH 1.4 ;
        PATH 54.0 22.3 54.0 25.5 ;
        WIDTH 1 ;
        PATH 54.5 3.3 54.5 26.0 ;
        WIDTH 0 ;
        PATH 44.0 10.8 44.0 9.3 25.3 9.3 ;
        WIDTH 1 ;
        PATH 25.5 9.5 43.0 9.5 43.0 11.5 43.8 11.5 ;
        WIDTH 1 ;
        PATH 42.0 21.8 42.0 16.0 38.5 16.0 38.5 12.8 38.3 12.8 ;
        
        LAYER ML1 ;
      # VIA 27 21.5 dcont
        RECT 26 20.5 28 22.5 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 33.5 21.5 dcont
        RECT 32.5 20.5 34.5 22.5 ;
      # VIA 27 23.5 dcont
        RECT 26 22.5 28 24.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 48 21.5 dcont
        RECT 47 20.5 49 22.5 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 38.5 23.5 dcont
        RECT 37.5 22.5 39.5 24.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 52 18.5 pcont
        RECT 51 17.5 53 19.5 ;
      # VIA 33.5 23.5 dcont
        RECT 32.5 22.5 34.5 24.5 ;
      # VIA 24 21.5 dcont
        RECT 23 20.5 25 22.5 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 40.5 6.5 pcont
        RECT 39.5 5.5 41.5 7.5 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 30.5 12 pcont
        RECT 29.5 11 31.5 13 ;
      # VIA 27.5 6.5 pcont
        RECT 26.5 5.5 28.5 7.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 49 16.5 pcont
        RECT 48 15.5 50 17.5 ;
      # VIA 39.5 3.5 dcont
        RECT 38.5 2.5 40.5 4.5 ;
      # VIA 28.5 18 pcont
        RECT 27.5 17 29.5 19 ;
      # VIA 33.5 25.5 dcont
        RECT 32.5 24.5 34.5 26.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 54 25.5 dcont
        RECT 53 24.5 55 26.5 ;
      # VIA 24 23.5 dcont
        RECT 23 22.5 25 24.5 ;
      # VIA 44.5 21.5 dcont
        RECT 43.5 20.5 45.5 22.5 ;
      # VIA 54 23.5 dcont
        RECT 53 22.5 55 24.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 27 25.5 dcont
        RECT 26 24.5 28 26.5 ;
      # VIA 54 21.5 dcont
        RECT 53 20.5 55 22.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 52 6.5 pcont
        RECT 51 5.5 53 7.5 ;
      # VIA 48 3.5 dcont
        RECT 47 2.5 49 4.5 ;
      # VIA 44.5 23.5 dcont
        RECT 43.5 22.5 45.5 24.5 ;
      # VIA 15 12 pcont
        RECT 14 11 16 13 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 25 10 pcont
        RECT 24 9 26 11 ;
      # VIA 31.5 15.5 pcont
        RECT 30.5 14.5 32.5 16.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 44.5 25.5 dcont
        RECT 43.5 24.5 45.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 38.5 21.5 dcont
        RECT 37.5 20.5 39.5 22.5 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 34.5 3.5 dcont
        RECT 33.5 2.5 35.5 4.5 ;
      # VIA 48 23.5 dcont
        RECT 47 22.5 49 24.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 29.5 3.5 dcont
        RECT 28.5 2.5 30.5 4.5 ;
      # VIA 38.5 25.5 dcont
        RECT 37.5 24.5 39.5 26.5 ;
      # VIA 54 3.5 dcont
        RECT 53 2.5 55 4.5 ;
      # VIA 20 6.5 pcont
        RECT 19 5.5 21 7.5 ;
      # VIA 35.5 13 pcont
        RECT 34.5 12 36.5 14 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 49 8.5 pcont
        RECT 48 7.5 50 9.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 44.5 3.5 dcont
        RECT 43.5 2.5 45.5 4.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 24 25.5 dcont
        RECT 23 24.5 25 26.5 ;
      # VIA 38.5 13 pcont
        RECT 37.5 12 39.5 14 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 41.5 21.5 dcont
        RECT 40.5 20.5 42.5 22.5 ;
      # VIA 48 25.5 dcont
        RECT 47 24.5 49 26.5 ;
      # VIA 41.5 25.5 dcont
        RECT 40.5 24.5 42.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 26 3.5 dcont
        RECT 25 2.5 27 4.5 ;
      # VIA 41.5 23.5 dcont
        RECT 40.5 22.5 42.5 24.5 ;
      # VIA 39.5 18.5 pcont
        RECT 38.5 17.5 40.5 19.5 ;
    END
END sff1
MACRO sff1_r
    CLASS core ;
    FOREIGN sff1_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 62.5 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN S
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.0 51.5 12.0 ;
        LAYER ML1 ;
        RECT 49.5 10.0 51.5 12.0 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 63.0 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 60.0 10.5 62.0 12.5 ;
        LAYER ML1 ;
        RECT 60.0 10.5 62.0 12.5 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 63.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 31.0 19.0 31.0 21.5 ;
        WIDTH 1 ;
        PATH 38.3 15.5 14.3 15.5 ;
        WIDTH 0 ;
        PATH 50.5 10.8 50.5 9.3 31.8 9.3 ;
        WIDTH 0 ;
        PATH 50.5 10.8 50.5 9.3 31.8 9.3 ;
        WIDTH 1 ;
        PATH 8.0 26.0 8.0 3.6 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 11.9 13.0 8.0 13.0 ;
        WIDTH 1 ;
        PATH 12.3 6.0 8.0 6.0 ;
        WIDTH 1 ;
        PATH 12.1 18.5 8.0 18.5 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        RECT 13.4 20.9 14.6 26.1 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 15.5 14.5 15.5 14.5 26.0 ;
        WIDTH 2 ;
        PATH 17.5 1.0 17.5 3.8 ;
        WIDTH 2 ;
        PATH 17.5 22.6 17.5 28.5 ;
        WIDTH 1 ;
        PATH 21.3 6.5 14.8 6.5 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 22.5 22.3 22.5 19.0 28.5 19.0 ;
        WIDTH 1 ;
        PATH 22.5 3.8 22.5 4.0 24.0 4.0 24.0 9.5 28.6 9.5 ;
        WIDTH 2 ;
        PATH 27.5 22.6 27.5 28.5 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.8 ;
        WIDTH 1 ;
        PATH 41.9 12.5 16.8 12.5 ;
        WIDTH 1 ;
        PATH 33.8 6.0 26.8 6.0 ;
        WIDTH 1.4 ;
        PATH 30.5 21.5 30.5 25.5 ;
        WIDTH 1 ;
        PATH 31.0 19.0 35.0 19.0 35.0 18.0 ;
        WIDTH 1 ;
        PATH 33.0 3.6 33.0 5.5 ;
        WIDTH 2 ;
        PATH 33.5 23.8 33.5 28.5 ;
        
        
        WIDTH 2 ;
        PATH 36.0 1.0 36.0 3.8 ;
        WIDTH 1.4 ;
        PATH 40.0 22.3 40.0 25.5 ;
        WIDTH 1 ;
        PATH 40.5 22.3 40.5 19.0 46.0 19.0 ;
        WIDTH 2 ;
        PATH 45.0 22.6 45.0 28.5 ;
        WIDTH 1 ;
        PATH 41.5 3.8 41.5 6.0 46.8 6.0 ;
        WIDTH 2 ;
        PATH 46.0 1.0 46.0 3.8 ;
        WIDTH 2 ;
        PATH 51.0 22.6 51.0 28.5 ;
        WIDTH 1 ;
        PATH 51.5 3.8 51.5 8.0 56.0 8.0 56.0 17.0 48.8 17.0 ;
        WIDTH 1.4 ;
        PATH 54.5 22.3 54.5 25.5 ;
        WIDTH 1 ;
        PATH 55.0 26.0 55.0 19.0 58.5 19.0 58.5 6.0 55.0 6.0 55.0 3.6 ;
        WIDTH 2 ;
        PATH 57.5 1.0 57.5 3.8 ;
        WIDTH 2 ;
        PATH 57.5 22.6 57.5 28.5 ;
        WIDTH 1.4 ;
        PATH 60.5 22.3 60.5 25.5 ;
        WIDTH 1 ;
        PATH 61.0 3.3 61.0 26.0 ;
        WIDTH 0 ;
        PATH 50.5 10.8 50.5 9.3 31.8 9.3 ;
        WIDTH 1 ;
        PATH 32.0 9.5 49.5 9.5 49.5 11.5 50.3 11.5 ;
        WIDTH 1 ;
        PATH 48.5 21.8 48.5 16.0 45.0 16.0 45.0 12.8 44.8 12.8 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        
        LAYER ML1 ;
      # VIA 5.5 13 pcont
        RECT 4.5 12 6.5 14 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 28.5 10 pcont
        RECT 27.5 9 29.5 11 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 40 21.5 dcont
        RECT 39 20.5 41 22.5 ;
      # VIA 33.5 23.5 dcont
        RECT 32.5 22.5 34.5 24.5 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 54.5 21.5 dcont
        RECT 53.5 20.5 55.5 22.5 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 45 23.5 dcont
        RECT 44 22.5 46 24.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 58.5 18.5 pcont
        RECT 57.5 17.5 59.5 19.5 ;
      # VIA 40 23.5 dcont
        RECT 39 22.5 41 24.5 ;
      # VIA 30.5 21.5 dcont
        RECT 29.5 20.5 31.5 22.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 47 6.5 pcont
        RECT 46 5.5 48 7.5 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 37 12 pcont
        RECT 36 11 38 13 ;
      # VIA 33.5 21.5 dcont
        RECT 32.5 20.5 34.5 22.5 ;
      # VIA 34 6.5 pcont
        RECT 33 5.5 35 7.5 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 55.5 16.5 pcont
        RECT 54.5 15.5 56.5 17.5 ;
      # VIA 46 3.5 dcont
        RECT 45 2.5 47 4.5 ;
      # VIA 35 18 pcont
        RECT 34 17 36 19 ;
      # VIA 40 25.5 dcont
        RECT 39 24.5 41 26.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 60.5 25.5 dcont
        RECT 59.5 24.5 61.5 26.5 ;
      # VIA 30.5 23.5 dcont
        RECT 29.5 22.5 31.5 24.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 60.5 23.5 dcont
        RECT 59.5 22.5 61.5 24.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 57.5 21.5 dcont
        RECT 56.5 20.5 58.5 22.5 ;
      # VIA 33.5 25.5 dcont
        RECT 32.5 24.5 34.5 26.5 ;
      # VIA 60.5 21.5 dcont
        RECT 59.5 20.5 61.5 22.5 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 58.5 6.5 pcont
        RECT 57.5 5.5 59.5 7.5 ;
      # VIA 54.5 3.5 dcont
        RECT 53.5 2.5 55.5 4.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 21.5 12 pcont
        RECT 20.5 11 22.5 13 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 31.5 10 pcont
        RECT 30.5 9 32.5 11 ;
      # VIA 38 15.5 pcont
        RECT 37 14.5 39 16.5 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 45 21.5 dcont
        RECT 44 20.5 46 22.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 57.5 23.5 dcont
        RECT 56.5 22.5 58.5 24.5 ;
      # VIA 41 3.5 dcont
        RECT 40 2.5 42 4.5 ;
      # VIA 54.5 23.5 dcont
        RECT 53.5 22.5 55.5 24.5 ;
      # VIA 57.5 25.5 dcont
        RECT 56.5 24.5 58.5 26.5 ;
      # VIA 36 3.5 dcont
        RECT 35 2.5 37 4.5 ;
      # VIA 45 25.5 dcont
        RECT 44 24.5 46 26.5 ;
      # VIA 60.5 3.5 dcont
        RECT 59.5 2.5 61.5 4.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 42 13 pcont
        RECT 41 12 43 14 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 55.5 8.5 pcont
        RECT 54.5 7.5 56.5 9.5 ;
      # VIA 57.5 3.5 dcont
        RECT 56.5 2.5 58.5 4.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 30.5 25.5 dcont
        RECT 29.5 24.5 31.5 26.5 ;
      # VIA 45 13 pcont
        RECT 44 12 46 14 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 48 21.5 dcont
        RECT 47 20.5 49 22.5 ;
      # VIA 54.5 25.5 dcont
        RECT 53.5 24.5 55.5 26.5 ;
      # VIA 48 25.5 dcont
        RECT 47 24.5 49 26.5 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 32.5 3.5 dcont
        RECT 31.5 2.5 33.5 4.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 48 23.5 dcont
        RECT 47 22.5 49 24.5 ;
      # VIA 46 18.5 pcont
        RECT 45 17.5 47 19.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
    END
END sff1_r
MACRO sff1m2
    CLASS core ;
    FOREIGN sff1m2 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 56.0 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
        RECT 3.5 9.0 5.5 11.0 ;
        LAYER ML1 ;
        RECT 3.5 9.0 5.5 11.0 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 53.5 10.5 55.5 12.5 ;
        LAYER ML1 ;
        RECT 53.5 10.5 55.5 12.5 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 11.0 9.0 13.0 11.0 ;
        LAYER ML1 ;
        RECT 11.0 9.0 13.0 11.0 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 56.5 30.0 ;
        END
    END VDD
    PIN S
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 43.0 10.5 45.0 12.5 ;
        LAYER ML1 ;
        RECT 43.0 10.5 45.0 12.5 ;
        END
    END S
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 56.5 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 24.5 19.0 24.5 21.4 ;
        WIDTH 1 ;
        PATH 1.5 26.0 1.5 3.6 ;
        WIDTH 1.4 ;
        PATH 1.5 22.3 1.5 25.5 ;
        WIDTH 1 ;
        PATH 5.3 13.0 1.8 13.0 ;
        WIDTH 1 ;
        PATH 5.6 18.5 1.5 18.5 ;
        WIDTH 1 ;
        PATH 5.9 6.0 1.5 6.0 ;
        WIDTH 2 ;
        PATH 4.5 22.6 4.5 28.5 ;
        WIDTH 2 ;
        PATH 4.5 1.0 4.5 3.8 ;
        WIDTH 1 ;
        PATH 8.0 3.6 8.0 9.5 7.5 9.5 7.5 16.0 8.0 16.0 8.0 26.0 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 1 ;
        PATH 15.0 6.0 8.0 6.0 ;
        WIDTH 1.4 ;
        PATH 16.0 22.3 16.0 25.5 ;
        WIDTH 1 ;
        PATH 16.0 22.3 16.0 18.5 22.0 18.5 ;
        WIDTH 1 ;
        PATH 16.3 3.8 16.3 4.0 17.5 4.0 17.5 10.0 22.4 10.0 ;
        WIDTH 1 ;
        PATH 8.3 16.0 31.3 16.0 ;
        WIDTH 2 ;
        PATH 21.0 22.6 21.0 28.5 ;
        WIDTH 2 ;
        PATH 21.0 1.0 21.0 3.8 ;
        WIDTH 1 ;
        PATH 33.5 13.0 10.3 13.0 ;
        WIDTH 1 ;
        PATH 26.4 6.0 20.5 6.0 ;
        WIDTH 1.4 ;
        PATH 24.0 21.5 24.0 25.5 ;
        WIDTH 1 ;
        PATH 24.5 19.0 27.8 19.0 27.8 18.7 ;
        WIDTH 1 ;
        PATH 26.5 3.5 26.5 6.1 ;
        WIDTH 2 ;
        PATH 27.0 23.8 27.0 28.5 ;
        
        
        WIDTH 2 ;
        PATH 29.5 1.0 29.5 3.8 ;
        WIDTH 1.4 ;
        PATH 32.0 22.3 32.0 25.5 ;
        WIDTH 1 ;
        PATH 25.6 10.0 44.5 10.0 ;
        WIDTH 1 ;
        PATH 32.5 22.6 32.5 19.0 38.5 19.0 ;
        WIDTH 2 ;
        PATH 37.0 22.6 37.0 28.5 ;
        WIDTH 1 ;
        PATH 35.0 3.8 35.0 6.0 40.3 6.0 ;
        WIDTH 2 ;
        PATH 39.5 1.0 39.5 3.8 ;
        WIDTH 1 ;
        PATH 40.5 14.0 40.5 21.5 ;
        WIDTH 2 ;
        PATH 43.0 22.6 43.0 28.5 ;
        WIDTH 1 ;
        PATH 45.0 3.8 45.0 8.0 48.5 8.0 48.5 14.0 38.4 14.0 ;
        WIDTH 1 ;
        PATH 49.3 17.0 40.5 17.0 ;
        WIDTH 1.4 ;
        PATH 48.0 22.3 48.0 25.5 ;
        WIDTH 1 ;
        PATH 48.5 26.0 48.5 19.0 52.0 19.0 52.0 6.0 48.5 6.0 48.5 3.6 ;
        WIDTH 2 ;
        PATH 51.0 1.0 51.0 3.8 ;
        WIDTH 2 ;
        PATH 51.0 22.6 51.0 28.5 ;
        WIDTH 1.4 ;
        PATH 54.0 22.3 54.0 25.5 ;
        WIDTH 1 ;
        PATH 54.5 3.3 54.5 26.0 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 22.5 18.7 22.5 10.0 ;
        WIDTH 1 ;
        PATH 28.0 18.4 28.0 6.0 ;
        WIDTH 1 ;
        PATH 38.0 18.7 38.0 7.0 41.0 7.0 ;
        LAYER ML1 ;
      # VIA 38 18.5 pcont
        RECT 37 17.5 39 19.5 ;
      # VIA 40 23.5 dcont
        RECT 39 22.5 41 24.5 ;
      # VIA 26 3.5 dcont
        RECT 25 2.5 27 4.5 ;
      # VIA 21 25.5 dcont
        RECT 20 24.5 22 26.5 ;
      # VIA 5.5 6.5 pcont
        RECT 4.5 5.5 6.5 7.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 40 25.5 dcont
        RECT 39 24.5 41 26.5 ;
      # VIA 48 25.5 dcont
        RECT 47 24.5 49 26.5 ;
      # VIA 40 21.5 dcont
        RECT 39 20.5 41 22.5 ;
      # VIA 16 21.5 dcont
        RECT 15 20.5 17 22.5 ;
      # VIA 16 3.5 dcont
        RECT 15 2.5 17 4.5 ;
      # VIA 7.5 3.5 dcont
        RECT 6.5 2.5 8.5 4.5 ;
      # VIA 38 14 pcont
        RECT 37 13 39 15 ;
      # VIA 24 25.5 dcont
        RECT 23 24.5 25 26.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 5.5 18.5 pcont
        RECT 4.5 17.5 6.5 19.5 ;
      # VIA 38 18.5 dcont
        RECT 37 17.5 39 19.5 ;
        LAYER ML2 ;
      # VIA 38 18.5 dcont
        RECT 37 17.5 39 19.5 ;
        LAYER ML1 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 44.5 3.5 dcont
        RECT 43.5 2.5 45.5 4.5 ;
      # VIA 16 23.5 dcont
        RECT 15 22.5 17 24.5 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML2 ;
      # VIA 22 10 dcont
        RECT 21 9 23 11 ;
        LAYER ML1 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 49 8.5 pcont
        RECT 48 7.5 50 9.5 ;
      # VIA 7.5 23.5 dcont
        RECT 6.5 22.5 8.5 24.5 ;
      # VIA 10 13 pcont
        RECT 9 12 11 14 ;
      # VIA 22 18.5 pcont
        RECT 21 17.5 23 19.5 ;
      # VIA 54 3.5 dcont
        RECT 53 2.5 55 4.5 ;
      # VIA 37 25.5 dcont
        RECT 36 24.5 38 26.5 ;
      # VIA 29.5 3.5 dcont
        RECT 28.5 2.5 30.5 4.5 ;
      # VIA 51 25.5 dcont
        RECT 50 24.5 52 26.5 ;
      # VIA 48 23.5 dcont
        RECT 47 22.5 49 24.5 ;
      # VIA 34.5 3.5 dcont
        RECT 33.5 2.5 35.5 4.5 ;
      # VIA 51 23.5 dcont
        RECT 50 22.5 52 24.5 ;
      # VIA 15 13 pcont
        RECT 14 12 16 14 ;
      # VIA 37 21.5 dcont
        RECT 36 20.5 38 22.5 ;
      # VIA 27 6.5 dcont
        RECT 26 5.5 28 7.5 ;
        LAYER ML2 ;
      # VIA 27 6.5 dcont
        RECT 26 5.5 28 7.5 ;
        LAYER ML1 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 16 25.5 dcont
        RECT 15 24.5 17 26.5 ;
      # VIA 43 25.5 dcont
        RECT 42 24.5 44 26.5 ;
      # VIA 5 13 pcont
        RECT 4 12 6 14 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 33 13.5 pcont
        RECT 32 12.5 34 14.5 ;
      # VIA 27 6.5 pcont
        RECT 26 5.5 28 7.5 ;
      # VIA 15 6.5 pcont
        RECT 14 5.5 16 7.5 ;
      # VIA 7.5 25.5 dcont
        RECT 6.5 24.5 8.5 26.5 ;
      # VIA 17 16 pcont
        RECT 16 15 18 17 ;
      # VIA 43 23.5 dcont
        RECT 42 22.5 44 24.5 ;
      # VIA 48 3.5 dcont
        RECT 47 2.5 49 4.5 ;
      # VIA 52 6.5 pcont
        RECT 51 5.5 53 7.5 ;
      # VIA 7.5 21.5 dcont
        RECT 6.5 20.5 8.5 22.5 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML2 ;
      # VIA 22 18.5 dcont
        RECT 21 17.5 23 19.5 ;
        LAYER ML1 ;
      # VIA 54 21.5 dcont
        RECT 53 20.5 55 22.5 ;
      # VIA 27 25.5 dcont
        RECT 26 24.5 28 26.5 ;
      # VIA 51 21.5 dcont
        RECT 50 20.5 52 22.5 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 21 21.5 dcont
        RECT 20 20.5 22 22.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 54 23.5 dcont
        RECT 53 22.5 55 24.5 ;
      # VIA 43 21.5 dcont
        RECT 42 20.5 44 22.5 ;
      # VIA 24 23.5 dcont
        RECT 23 22.5 25 24.5 ;
      # VIA 54 25.5 dcont
        RECT 53 24.5 55 26.5 ;
      # VIA 21 23.5 dcont
        RECT 20 22.5 22 24.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
      # VIA 32 25.5 dcont
        RECT 31 24.5 33 26.5 ;
      # VIA 28 13 pcont
        RECT 27 12 29 14 ;
      # VIA 39.5 3.5 dcont
        RECT 38.5 2.5 40.5 4.5 ;
      # VIA 28 18.5 dcont
        RECT 27 17.5 29 19.5 ;
        LAYER ML2 ;
      # VIA 28 18.5 dcont
        RECT 27 17.5 29 19.5 ;
        LAYER ML1 ;
      # VIA 49 16.5 pcont
        RECT 48 15.5 50 17.5 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 28 18.5 pcont
        RECT 27 17.5 29 19.5 ;
      # VIA 31 16.5 pcont
        RECT 30 15.5 32 17.5 ;
      # VIA 40.5 6.5 dcont
        RECT 39.5 5.5 41.5 7.5 ;
        LAYER ML2 ;
      # VIA 40.5 6.5 dcont
        RECT 39.5 5.5 41.5 7.5 ;
        LAYER ML1 ;
      # VIA 40.5 6.5 pcont
        RECT 39.5 5.5 41.5 7.5 ;
      # VIA 20 6.5 pcont
        RECT 19 5.5 21 7.5 ;
      # VIA 24 21.5 dcont
        RECT 23 20.5 25 22.5 ;
      # VIA 32 23.5 dcont
        RECT 31 22.5 33 24.5 ;
      # VIA 52 18.5 pcont
        RECT 51 17.5 53 19.5 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 37 23.5 dcont
        RECT 36 22.5 38 24.5 ;
      # VIA 21 3.5 dcont
        RECT 20 2.5 22 4.5 ;
      # VIA 22 10 pcont
        RECT 21 9 23 11 ;
      # VIA 48 21.5 dcont
        RECT 47 20.5 49 22.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 27 23.5 dcont
        RECT 26 22.5 28 24.5 ;
      # VIA 32 21.5 dcont
        RECT 31 20.5 33 22.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 25.5 10 pcont
        RECT 24.5 9 26.5 11 ;
      # VIA 27 21.5 dcont
        RECT 26 20.5 28 22.5 ;
    END
END sff1m2
MACRO sff1m2_r
    CLASS core ;
    FOREIGN sff1m2_r 0.0 0.0 ;
    ORIGIN 0.0 0.0 ;
    SIZE 62.5 BY 29.0 ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER ML2 ;
         RECT 1.0 14.5 3.0 16.5 ;
        LAYER ML1 ;
        RECT 1.0 14.5 3.0 16.5 ;
        END
    END CK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.5 28.0 63.0 30.0 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 17.5 9.0 19.5 11.0 ;
        LAYER ML1 ;
        RECT 17.5 9.0 19.5 11.0 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 60.0 10.5 62.0 12.5 ;
        LAYER ML1 ;
        RECT 60.0 10.5 62.0 12.5 ;
        END
    END Q
    PIN S
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 49.5 10.5 51.5 12.5 ;
        LAYER ML1 ;
        RECT 49.5 10.5 51.5 12.5 ;
        END
    END S
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.5 -1.0 63.0 1.0 ;
        END
    END VSS
    OBS
        LAYER ML1 ;
        
        WIDTH 1 ;
        PATH 31.0 19.0 31.0 21.4 ;
        WIDTH 1 ;
        PATH 8.0 26.0 8.0 3.6 ;
        WIDTH 1.4 ;
        PATH 8.0 22.3 8.0 25.5 ;
        WIDTH 1 ;
        PATH 11.8 13.0 8.3 13.0 ;
        WIDTH 1 ;
        PATH 12.1 18.5 8.0 18.5 ;
        WIDTH 1 ;
        PATH 12.4 6.0 8.0 6.0 ;
        WIDTH 2 ;
        PATH 11.0 22.6 11.0 28.5 ;
        WIDTH 2 ;
        PATH 11.0 1.0 11.0 3.8 ;
        WIDTH 1 ;
        PATH 14.5 3.6 14.5 9.5 14.0 9.5 14.0 16.0 14.5 16.0 14.5 26.0 ;
        WIDTH 2 ;
        PATH 17.5 1.0 17.5 3.8 ;
        WIDTH 2 ;
        PATH 17.5 22.6 17.5 28.5 ;
        WIDTH 1 ;
        PATH 21.5 6.0 14.5 6.0 ;
        WIDTH 1.4 ;
        PATH 22.5 22.3 22.5 25.5 ;
        WIDTH 1 ;
        PATH 22.5 22.3 22.5 18.5 28.5 18.5 ;
        WIDTH 1 ;
        PATH 22.8 3.8 22.8 4.0 24.0 4.0 24.0 10.0 28.9 10.0 ;
        WIDTH 1 ;
        PATH 14.8 16.0 37.8 16.0 ;
        WIDTH 2 ;
        PATH 27.5 22.6 27.5 28.5 ;
        WIDTH 2 ;
        PATH 27.5 1.0 27.5 3.8 ;
        WIDTH 1 ;
        PATH 40.0 13.0 16.8 13.0 ;
        WIDTH 1 ;
        PATH 32.9 6.0 27.0 6.0 ;
        WIDTH 1.4 ;
        PATH 30.5 21.5 30.5 25.5 ;
        WIDTH 1 ;
        PATH 31.0 19.0 34.3 19.0 34.3 18.7 ;
        WIDTH 1 ;
        PATH 33.0 3.5 33.0 6.1 ;
        WIDTH 2 ;
        PATH 33.5 23.8 33.5 28.5 ;
        
        
        WIDTH 2 ;
        PATH 36.0 1.0 36.0 3.8 ;
        WIDTH 1.4 ;
        PATH 38.5 22.3 38.5 25.5 ;
        WIDTH 1 ;
        PATH 32.1 10.0 51.0 10.0 ;
        WIDTH 1 ;
        PATH 39.0 22.6 39.0 19.0 45.0 19.0 ;
        WIDTH 2 ;
        PATH 43.5 22.6 43.5 28.5 ;
        WIDTH 1 ;
        PATH 41.5 3.8 41.5 6.0 46.8 6.0 ;
        WIDTH 2 ;
        PATH 46.0 1.0 46.0 3.8 ;
        WIDTH 1 ;
        PATH 47.0 14.0 47.0 21.5 ;
        WIDTH 2 ;
        PATH 49.5 22.6 49.5 28.5 ;
        WIDTH 1 ;
        PATH 51.5 3.8 51.5 8.0 55.0 8.0 55.0 14.0 44.9 14.0 ;
        WIDTH 1 ;
        PATH 55.8 17.0 47.0 17.0 ;
        WIDTH 1.4 ;
        PATH 54.5 22.3 54.5 25.5 ;
        WIDTH 1 ;
        PATH 55.0 26.0 55.0 19.0 58.5 19.0 58.5 6.0 55.0 6.0 55.0 3.6 ;
        WIDTH 2 ;
        PATH 57.5 1.0 57.5 3.8 ;
        WIDTH 2 ;
        PATH 57.5 22.6 57.5 28.5 ;
        WIDTH 1.4 ;
        PATH 60.5 22.3 60.5 25.5 ;
        WIDTH 1 ;
        PATH 61.0 3.3 61.0 26.0 ;
        WIDTH 2 ;
        PATH 1.5 21.5 1.5 28.5 ;
        WIDTH 2 ;
        PATH 1.5 1.0 1.5 3.5 ;
        
        
        WIDTH 1.4 ;
        PATH 4.5 22.3 4.5 25.5 ;
        WIDTH 1 ;
        PATH 4.5 20.5 4.5 3.8 ;
        
       LAYER ML2 ;
        WIDTH 1 ;
        PATH 29.0 18.7 29.0 10.0 ;
        WIDTH 1 ;
        PATH 34.5 18.4 34.5 6.0 ;
        WIDTH 1 ;
        PATH 44.5 18.7 44.5 7.0 47.5 7.0 ;
        LAYER ML1 ;
      # VIA 5.5 13 pcont
        RECT 4.5 12 6.5 14 ;
      # VIA 1.5 21.5 dcont
        RECT 0.5 20.5 2.5 22.5 ;
      # VIA 1.5 3.5 dcont
        RECT 0.5 2.5 2.5 4.5 ;
      # VIA 1.5 25.5 dcont
        RECT 0.5 24.5 2.5 26.5 ;
      # VIA 4.5 23.5 dcont
        RECT 3.5 22.5 5.5 24.5 ;
      # VIA 44.5 18.5 pcont
        RECT 43.5 17.5 45.5 19.5 ;
      # VIA 46.5 23.5 dcont
        RECT 45.5 22.5 47.5 24.5 ;
      # VIA 32.5 3.5 dcont
        RECT 31.5 2.5 33.5 4.5 ;
      # VIA 27.5 25.5 dcont
        RECT 26.5 24.5 28.5 26.5 ;
      # VIA 12 6.5 pcont
        RECT 11 5.5 13 7.5 ;
      # VIA 8 23.5 dcont
        RECT 7 22.5 9 24.5 ;
      # VIA 46.5 25.5 dcont
        RECT 45.5 24.5 47.5 26.5 ;
      # VIA 54.5 25.5 dcont
        RECT 53.5 24.5 55.5 26.5 ;
      # VIA 46.5 21.5 dcont
        RECT 45.5 20.5 47.5 22.5 ;
      # VIA 22.5 21.5 dcont
        RECT 21.5 20.5 23.5 22.5 ;
      # VIA 22.5 3.5 dcont
        RECT 21.5 2.5 23.5 4.5 ;
      # VIA 14 3.5 dcont
        RECT 13 2.5 15 4.5 ;
      # VIA 44.5 14 pcont
        RECT 43.5 13 45.5 15 ;
      # VIA 30.5 25.5 dcont
        RECT 29.5 24.5 31.5 26.5 ;
      # VIA 8 3.5 dcont
        RECT 7 2.5 9 4.5 ;
      # VIA 44.5 18.5 dcont
        RECT 43.5 17.5 45.5 19.5 ;
        LAYER ML2 ;
      # VIA 44.5 18.5 dcont
        RECT 43.5 17.5 45.5 19.5 ;
        LAYER ML1 ;
      # VIA 12 18.5 pcont
        RECT 11 17.5 13 19.5 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML2 ;
      # VIA 28.5 10 dcont
        RECT 27.5 9 29.5 11 ;
        LAYER ML1 ;
      # VIA 11 3.5 dcont
        RECT 10 2.5 12 4.5 ;
      # VIA 51 3.5 dcont
        RECT 50 2.5 52 4.5 ;
      # VIA 22.5 23.5 dcont
        RECT 21.5 22.5 23.5 24.5 ;
      # VIA 57.5 3.5 dcont
        RECT 56.5 2.5 58.5 4.5 ;
      # VIA 55.5 8.5 pcont
        RECT 54.5 7.5 56.5 9.5 ;
      # VIA 14 23.5 dcont
        RECT 13 22.5 15 24.5 ;
      # VIA 16.5 13 pcont
        RECT 15.5 12 17.5 14 ;
      # VIA 28.5 18.5 pcont
        RECT 27.5 17.5 29.5 19.5 ;
      # VIA 60.5 3.5 dcont
        RECT 59.5 2.5 61.5 4.5 ;
      # VIA 43.5 25.5 dcont
        RECT 42.5 24.5 44.5 26.5 ;
      # VIA 36 3.5 dcont
        RECT 35 2.5 37 4.5 ;
      # VIA 57.5 25.5 dcont
        RECT 56.5 24.5 58.5 26.5 ;
      # VIA 54.5 23.5 dcont
        RECT 53.5 22.5 55.5 24.5 ;
      # VIA 41 3.5 dcont
        RECT 40 2.5 42 4.5 ;
      # VIA 57.5 23.5 dcont
        RECT 56.5 22.5 58.5 24.5 ;
      # VIA 21.5 13 pcont
        RECT 20.5 12 22.5 14 ;
      # VIA 43.5 21.5 dcont
        RECT 42.5 20.5 44.5 22.5 ;
      # VIA 33.5 6.5 dcont
        RECT 32.5 5.5 34.5 7.5 ;
        LAYER ML2 ;
      # VIA 33.5 6.5 dcont
        RECT 32.5 5.5 34.5 7.5 ;
        LAYER ML1 ;
      # VIA 11 25.5 dcont
        RECT 10 24.5 12 26.5 ;
      # VIA 22.5 25.5 dcont
        RECT 21.5 24.5 23.5 26.5 ;
      # VIA 49.5 25.5 dcont
        RECT 48.5 24.5 50.5 26.5 ;
      # VIA 11.5 13 pcont
        RECT 10.5 12 12.5 14 ;
      # VIA 17.5 21.5 dcont
        RECT 16.5 20.5 18.5 22.5 ;
      # VIA 39.5 13.5 pcont
        RECT 38.5 12.5 40.5 14.5 ;
      # VIA 33.5 6.5 pcont
        RECT 32.5 5.5 34.5 7.5 ;
      # VIA 21.5 6.5 pcont
        RECT 20.5 5.5 22.5 7.5 ;
      # VIA 14 25.5 dcont
        RECT 13 24.5 15 26.5 ;
      # VIA 23.5 16 pcont
        RECT 22.5 15 24.5 17 ;
      # VIA 49.5 23.5 dcont
        RECT 48.5 22.5 50.5 24.5 ;
      # VIA 54.5 3.5 dcont
        RECT 53.5 2.5 55.5 4.5 ;
      # VIA 33.5 21.5 dcont
        RECT 32.5 20.5 34.5 22.5 ;
      # VIA 58.5 6.5 pcont
        RECT 57.5 5.5 59.5 7.5 ;
      # VIA 14 21.5 dcont
        RECT 13 20.5 15 22.5 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML2 ;
      # VIA 28.5 18.5 dcont
        RECT 27.5 17.5 29.5 19.5 ;
        LAYER ML1 ;
      # VIA 60.5 21.5 dcont
        RECT 59.5 20.5 61.5 22.5 ;
      # VIA 33.5 25.5 dcont
        RECT 32.5 24.5 34.5 26.5 ;
      # VIA 57.5 21.5 dcont
        RECT 56.5 20.5 58.5 22.5 ;
      # VIA 17.5 3.5 dcont
        RECT 16.5 2.5 18.5 4.5 ;
      # VIA 27.5 21.5 dcont
        RECT 26.5 20.5 28.5 22.5 ;
      # VIA 11 23.5 dcont
        RECT 10 22.5 12 24.5 ;
      # VIA 60.5 23.5 dcont
        RECT 59.5 22.5 61.5 24.5 ;
      # VIA 49.5 21.5 dcont
        RECT 48.5 20.5 50.5 22.5 ;
      # VIA 30.5 23.5 dcont
        RECT 29.5 22.5 31.5 24.5 ;
      # VIA 60.5 25.5 dcont
        RECT 59.5 24.5 61.5 26.5 ;
      # VIA 27.5 23.5 dcont
        RECT 26.5 22.5 28.5 24.5 ;
      # VIA 11 21.5 dcont
        RECT 10 20.5 12 22.5 ;
      # VIA 38.5 25.5 dcont
        RECT 37.5 24.5 39.5 26.5 ;
      # VIA 34.5 13 pcont
        RECT 33.5 12 35.5 14 ;
      # VIA 46 3.5 dcont
        RECT 45 2.5 47 4.5 ;
      # VIA 34.5 18.5 dcont
        RECT 33.5 17.5 35.5 19.5 ;
        LAYER ML2 ;
      # VIA 34.5 18.5 dcont
        RECT 33.5 17.5 35.5 19.5 ;
        LAYER ML1 ;
      # VIA 55.5 16.5 pcont
        RECT 54.5 15.5 56.5 17.5 ;
      # VIA 17.5 25.5 dcont
        RECT 16.5 24.5 18.5 26.5 ;
      # VIA 34.5 18.5 pcont
        RECT 33.5 17.5 35.5 19.5 ;
      # VIA 47 6.5 dcont
        RECT 46 5.5 48 7.5 ;
        LAYER ML2 ;
      # VIA 47 6.5 dcont
        RECT 46 5.5 48 7.5 ;
        LAYER ML1 ;
      # VIA 37.5 16.5 pcont
        RECT 36.5 15.5 38.5 17.5 ;
      # VIA 47 6.5 pcont
        RECT 46 5.5 48 7.5 ;
      # VIA 26.5 6.5 pcont
        RECT 25.5 5.5 27.5 7.5 ;
      # VIA 30.5 21.5 dcont
        RECT 29.5 20.5 31.5 22.5 ;
      # VIA 38.5 23.5 dcont
        RECT 37.5 22.5 39.5 24.5 ;
      # VIA 58.5 18.5 pcont
        RECT 57.5 17.5 59.5 19.5 ;
      # VIA 8 21.5 dcont
        RECT 7 20.5 9 22.5 ;
      # VIA 43.5 23.5 dcont
        RECT 42.5 22.5 44.5 24.5 ;
      # VIA 27.5 3.5 dcont
        RECT 26.5 2.5 28.5 4.5 ;
      # VIA 28.5 10 pcont
        RECT 27.5 9 29.5 11 ;
      # VIA 54.5 21.5 dcont
        RECT 53.5 20.5 55.5 22.5 ;
      # VIA 17.5 23.5 dcont
        RECT 16.5 22.5 18.5 24.5 ;
      # VIA 33.5 23.5 dcont
        RECT 32.5 22.5 34.5 24.5 ;
      # VIA 38.5 21.5 dcont
        RECT 37.5 20.5 39.5 22.5 ;
      # VIA 8 25.5 dcont
        RECT 7 24.5 9 26.5 ;
      # VIA 32 10 pcont
        RECT 31 9 33 11 ;
      # VIA 4.5 25.5 dcont
        RECT 3.5 24.5 5.5 26.5 ;
      # VIA 1.5 23.5 dcont
        RECT 0.5 22.5 2.5 24.5 ;
      # VIA 4.5 3.5 dcont
        RECT 3.5 2.5 5.5 4.5 ;
      # VIA 4.5 21.5 dcont
        RECT 3.5 20.5 5.5 22.5 ;
    END
END sff1m2_r


END LIBRARY
