# C:/Users/akita/Documents/or31.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:43:39 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO or31
    CLASS core ;
    FOREIGN or31 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 18.500 BY 32.500 ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 16.000 30.000 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.000 11.500 6.000 13.500 ;
        LAYER ML1 ;
        RECT 4.000 11.500 6.000 13.500 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.000 9.000 15.000 11.000 ;
        LAYER ML1 ;
        RECT 13.000 9.000 15.000 11.000 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.000 12.000 9.000 14.000 ;
        LAYER ML1 ;
        RECT 7.000 12.000 9.000 14.000 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 16.000 1.000 ;
        END
    END VSS
    OBS
    END
END or31

END LIBRARY
