# C:/Users/akita/Documents/sff1_r.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:44:54 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO sff1_r
    CLASS core ;
    FOREIGN sff1_r -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 65.500 BY 32.500 ;
    PIN CK
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END CK
    PIN S
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER ML2 ;
        RECT 49.500 10.000 51.500 12.000 ;
        LAYER ML1 ;
        RECT 49.500 10.000 51.500 12.000 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 63.000 30.000 ;
        END
    END VDD
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 17.500 9.000 19.500 11.000 ;
        LAYER ML1 ;
        RECT 17.500 9.000 19.500 11.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 60.000 10.500 62.000 12.500 ;
        LAYER ML1 ;
        RECT 60.000 10.500 62.000 12.500 ;
        END
    END Q
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 63.000 1.000 ;
        END
    END VSS
    OBS
    END
END sff1_r

END LIBRARY
