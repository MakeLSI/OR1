# C:/Users/akita/Documents/or21.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:43:29 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO or21
    CLASS core ;
    FOREIGN or21 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 15.500 BY 32.500 ;
    PIN 
        DIRECTION INPUT ;
        USE POWER ;
        END
    END 
    PIN Y
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.000 8.000 12.000 10.000 ;
        LAYER ML1 ;
        RECT 10.000 8.000 12.000 10.000 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 13.000 30.000 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.000 11.500 6.000 13.500 ;
        LAYER ML1 ;
        RECT 4.000 11.500 6.000 13.500 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 8.500 3.000 10.500 ;
        LAYER ML1 ;
        RECT 1.000 8.500 3.000 10.500 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 13.000 1.000 ;
        END
    END VSS
    OBS
    END
END or21

END LIBRARY
