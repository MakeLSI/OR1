# C:/Users/akita/Documents/na222.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:37:09 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO na222
    CLASS core ;
    FOREIGN na222 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 18.500 BY 32.500 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.000 10.500 15.000 12.500 ;
        LAYER ML1 ;
        RECT 13.000 10.500 15.000 12.500 ;
        END
    END YB
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.000 10.000 6.000 12.000 ;
        LAYER ML1 ;
        RECT 4.000 10.000 6.000 12.000 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 16.000 30.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 16.000 1.000 ;
        END
    END VSS
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.000 14.500 12.000 16.500 ;
        LAYER ML1 ;
        RECT 10.000 14.500 12.000 16.500 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.000 11.500 9.000 13.500 ;
        LAYER ML1 ;
        RECT 7.000 11.500 9.000 13.500 ;
        END
    END B1
    OBS
    END
END na222

END LIBRARY
