# C:/Users/akita/Documents/exnr.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:35:17 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO exnr
    CLASS core ;
    FOREIGN exnr -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 25.000 BY 32.500 ;
    PIN 
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT 23.500 7.000 23.500 7.000 ;
        END
    END 
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 3.000 10.500 5.000 12.500 ;
        LAYER ML1 ;
        RECT 3.000 10.500 5.000 12.500 ;
        END
    END B
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 21.500 30.000 ;
        END
    END VDD
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 18.500 12.500 20.500 14.500 ;
        LAYER ML1 ;
        RECT 18.500 12.500 20.500 14.500 ;
        END
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 21.500 1.000 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 6.000 13.500 8.000 15.500 ;
        LAYER ML1 ;
        RECT 6.000 13.500 8.000 15.500 ;
        END
    END A
    OBS
    END
END exnr

END LIBRARY
