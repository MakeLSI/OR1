# C:/Users/akita/Documents/inv1lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:35:41 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO inv1
    CLASS core ;
    FOREIGN inv1 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 9.500 BY 32.500 ;
    PIN 
        DIRECTION INPUT ;
        USE POWER ;
        END
    END 
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.000 10.500 6.000 12.500 ;
        END
    END YB
    PIN X
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 4.000 10.500 6.000 12.500 ;
        END
    END X
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 7.000 30.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER FRAME ;
        RECT -0.500 -1.000 7.000 1.000 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END A
    OBS
    END
END inv1

END LIBRARY
