# C:/Users/akita/Documents/ttt.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:32:22 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO buf2
    CLASS core ;
    FOREIGN buf2 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 15.500 BY 32.500 ;
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.000 14.000 9.000 16.000 ;
        LAYER ML1 ;
        RECT 7.000 14.000 9.000 16.000 ;
        END
    END Y
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 13.000 30.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 13.000 1.000 ;
        END
    END VSS
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END A
    OBS
    END
END buf2

END LIBRARY
