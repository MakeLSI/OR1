# C:/Users/akita/Documents/sff1m2.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:45:04 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO sff1m2
    CLASS core ;
    FOREIGN sff1m2 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 59.000 BY 32.500 ;
    PIN CK
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 3.500 9.000 5.500 11.000 ;
        LAYER ML1 ;
        RECT 3.500 9.000 5.500 11.000 ;
        END
    END CK
    PIN Q
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 53.500 10.500 55.500 12.500 ;
        LAYER ML1 ;
        RECT 53.500 10.500 55.500 12.500 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 11.000 9.000 13.000 11.000 ;
        LAYER ML1 ;
        RECT 11.000 9.000 13.000 11.000 ;
        END
    END D
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 56.500 30.000 ;
        END
    END VDD
    PIN S
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER ML2 ;
        RECT 43.000 10.500 45.000 12.500 ;
        LAYER ML1 ;
        RECT 43.000 10.500 45.000 12.500 ;
        END
    END S
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 56.500 1.000 ;
        END
    END VSS
    OBS
    END
END sff1m2

END LIBRARY
