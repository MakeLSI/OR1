# C:/Users/akita/Documents/na212.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:36:59 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO na212
    CLASS core ;
    FOREIGN na212 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 15.500 BY 32.500 ;
    PIN 
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER FRAME ;
        RECT 12.000 12.500 13.000 12.500 ;
        END
    END 
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 10.000 8.500 12.000 10.500 ;
        LAYER ML1 ;
        RECT 10.000 8.500 12.000 10.500 ;
        END
    END YB
    PIN A1
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 4.000 11.500 6.000 13.500 ;
        RECT 4.000 11.500 6.000 13.500 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END A0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 13.000 30.000 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 13.000 1.000 ;
        END
    END VSS
    PIN B0
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML1 ;
        RECT 7.000 12.000 9.000 14.000 ;
        RECT 7.000 12.000 9.000 14.000 ;
        END
    END B0
    OBS
    END
END na212

END LIBRARY
