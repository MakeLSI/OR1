# C:/Users/akita/Documents/na41.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:37:29 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO na41
    CLASS core ;
    FOREIGN na41 -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 18.500 BY 32.500 ;
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 13.000 9.500 15.000 11.500 ;
        LAYER ML1 ;
        RECT 13.000 9.500 15.000 11.500 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 16.000 30.000 ;
        END
    END VDD
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 4.000 12.500 6.000 14.500 ;
        LAYER ML1 ;
        RECT 4.000 12.500 6.000 14.500 ;
        END
    END B
    PIN D
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER ML2 ;
        RECT 10.000 6.500 12.000 8.500 ;
        LAYER ML1 ;
        RECT 10.000 6.500 12.000 8.500 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 7.000 9.500 9.000 11.500 ;
        LAYER ML1 ;
        RECT 7.000 9.500 9.000 11.500 ;
        END
    END C
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 15.500 3.000 17.500 ;
        LAYER ML1 ;
        RECT 1.000 15.500 3.000 17.500 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 16.000 1.000 ;
        END
    END VSS
    OBS
    END
END na41

END LIBRARY
