# C:/Users/akita/Documents/000.lef
# Created by Glade release version 4.7.35 compiled on May 19 2020 19:14:35
# Run by akita on host LAPTOP-E0CJ65QR at Wed Jun  3 17:33:17 2020

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO cinv
    CLASS core ;
    FOREIGN cinv -1.500 -1.500 ;
    ORIGIN 1.500 1.500 ;
    SIZE 14.500 BY 32.500 ;
    PIN OE
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 1.000 14.500 3.000 16.500 ;
        LAYER ML1 ;
        RECT 1.000 14.500 3.000 16.500 ;
        END
    END OE
    PIN YB
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 9.000 7.500 11.000 9.500 ;
        LAYER ML1 ;
        RECT 9.000 7.500 11.000 9.500 ;
        END
    END YB
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        PORT
        LAYER ML1 ;
        RECT -0.500 28.000 12.000 30.000 ;
        END
    END VDD
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER ML2 ;
        RECT 6.500 11.500 8.500 13.500 ;
        LAYER ML1 ;
        RECT 6.500 11.500 8.500 13.500 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        PORT
        LAYER ML1 ;
        RECT -0.500 -1.000 12.000 1.000 ;
        END
    END VSS
    OBS
    END
END cinv

END LIBRARY
